module STORE_QUEUE_LSQ_a( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_bbStart, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_0, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_1, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_2, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_3, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_4, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_5, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_6, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_7, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_8, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_9, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_10, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_11, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_12, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_13, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_14, // @[:@6.4]
  input  [3:0]  io_bbStoreOffsets_15, // @[:@6.4]
  input         io_bbNumStores, // @[:@6.4]
  output [3:0]  io_storeTail, // @[:@6.4]
  output [3:0]  io_storeHead, // @[:@6.4]
  output        io_storeEmpty, // @[:@6.4]
  input  [3:0]  io_loadTail, // @[:@6.4]
  input  [3:0]  io_loadHead, // @[:@6.4]
  input         io_loadEmpty, // @[:@6.4]
  input         io_loadAddressDone_0, // @[:@6.4]
  input         io_loadAddressDone_1, // @[:@6.4]
  input         io_loadAddressDone_2, // @[:@6.4]
  input         io_loadAddressDone_3, // @[:@6.4]
  input         io_loadAddressDone_4, // @[:@6.4]
  input         io_loadAddressDone_5, // @[:@6.4]
  input         io_loadAddressDone_6, // @[:@6.4]
  input         io_loadAddressDone_7, // @[:@6.4]
  input         io_loadAddressDone_8, // @[:@6.4]
  input         io_loadAddressDone_9, // @[:@6.4]
  input         io_loadAddressDone_10, // @[:@6.4]
  input         io_loadAddressDone_11, // @[:@6.4]
  input         io_loadAddressDone_12, // @[:@6.4]
  input         io_loadAddressDone_13, // @[:@6.4]
  input         io_loadAddressDone_14, // @[:@6.4]
  input         io_loadAddressDone_15, // @[:@6.4]
  input         io_loadDataDone_0, // @[:@6.4]
  input         io_loadDataDone_1, // @[:@6.4]
  input         io_loadDataDone_2, // @[:@6.4]
  input         io_loadDataDone_3, // @[:@6.4]
  input         io_loadDataDone_4, // @[:@6.4]
  input         io_loadDataDone_5, // @[:@6.4]
  input         io_loadDataDone_6, // @[:@6.4]
  input         io_loadDataDone_7, // @[:@6.4]
  input         io_loadDataDone_8, // @[:@6.4]
  input         io_loadDataDone_9, // @[:@6.4]
  input         io_loadDataDone_10, // @[:@6.4]
  input         io_loadDataDone_11, // @[:@6.4]
  input         io_loadDataDone_12, // @[:@6.4]
  input         io_loadDataDone_13, // @[:@6.4]
  input         io_loadDataDone_14, // @[:@6.4]
  input         io_loadDataDone_15, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_0, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_1, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_2, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_3, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_4, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_5, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_6, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_7, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_8, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_9, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_10, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_11, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_12, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_13, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_14, // @[:@6.4]
  input  [30:0] io_loadAddressQueue_15, // @[:@6.4]
  output        io_storeAddrDone_0, // @[:@6.4]
  output        io_storeAddrDone_1, // @[:@6.4]
  output        io_storeAddrDone_2, // @[:@6.4]
  output        io_storeAddrDone_3, // @[:@6.4]
  output        io_storeAddrDone_4, // @[:@6.4]
  output        io_storeAddrDone_5, // @[:@6.4]
  output        io_storeAddrDone_6, // @[:@6.4]
  output        io_storeAddrDone_7, // @[:@6.4]
  output        io_storeAddrDone_8, // @[:@6.4]
  output        io_storeAddrDone_9, // @[:@6.4]
  output        io_storeAddrDone_10, // @[:@6.4]
  output        io_storeAddrDone_11, // @[:@6.4]
  output        io_storeAddrDone_12, // @[:@6.4]
  output        io_storeAddrDone_13, // @[:@6.4]
  output        io_storeAddrDone_14, // @[:@6.4]
  output        io_storeAddrDone_15, // @[:@6.4]
  output        io_storeDataDone_0, // @[:@6.4]
  output        io_storeDataDone_1, // @[:@6.4]
  output        io_storeDataDone_2, // @[:@6.4]
  output        io_storeDataDone_3, // @[:@6.4]
  output        io_storeDataDone_4, // @[:@6.4]
  output        io_storeDataDone_5, // @[:@6.4]
  output        io_storeDataDone_6, // @[:@6.4]
  output        io_storeDataDone_7, // @[:@6.4]
  output        io_storeDataDone_8, // @[:@6.4]
  output        io_storeDataDone_9, // @[:@6.4]
  output        io_storeDataDone_10, // @[:@6.4]
  output        io_storeDataDone_11, // @[:@6.4]
  output        io_storeDataDone_12, // @[:@6.4]
  output        io_storeDataDone_13, // @[:@6.4]
  output        io_storeDataDone_14, // @[:@6.4]
  output        io_storeDataDone_15, // @[:@6.4]
  output [30:0] io_storeAddrQueue_0, // @[:@6.4]
  output [30:0] io_storeAddrQueue_1, // @[:@6.4]
  output [30:0] io_storeAddrQueue_2, // @[:@6.4]
  output [30:0] io_storeAddrQueue_3, // @[:@6.4]
  output [30:0] io_storeAddrQueue_4, // @[:@6.4]
  output [30:0] io_storeAddrQueue_5, // @[:@6.4]
  output [30:0] io_storeAddrQueue_6, // @[:@6.4]
  output [30:0] io_storeAddrQueue_7, // @[:@6.4]
  output [30:0] io_storeAddrQueue_8, // @[:@6.4]
  output [30:0] io_storeAddrQueue_9, // @[:@6.4]
  output [30:0] io_storeAddrQueue_10, // @[:@6.4]
  output [30:0] io_storeAddrQueue_11, // @[:@6.4]
  output [30:0] io_storeAddrQueue_12, // @[:@6.4]
  output [30:0] io_storeAddrQueue_13, // @[:@6.4]
  output [30:0] io_storeAddrQueue_14, // @[:@6.4]
  output [30:0] io_storeAddrQueue_15, // @[:@6.4]
  output [31:0] io_storeDataQueue_0, // @[:@6.4]
  output [31:0] io_storeDataQueue_1, // @[:@6.4]
  output [31:0] io_storeDataQueue_2, // @[:@6.4]
  output [31:0] io_storeDataQueue_3, // @[:@6.4]
  output [31:0] io_storeDataQueue_4, // @[:@6.4]
  output [31:0] io_storeDataQueue_5, // @[:@6.4]
  output [31:0] io_storeDataQueue_6, // @[:@6.4]
  output [31:0] io_storeDataQueue_7, // @[:@6.4]
  output [31:0] io_storeDataQueue_8, // @[:@6.4]
  output [31:0] io_storeDataQueue_9, // @[:@6.4]
  output [31:0] io_storeDataQueue_10, // @[:@6.4]
  output [31:0] io_storeDataQueue_11, // @[:@6.4]
  output [31:0] io_storeDataQueue_12, // @[:@6.4]
  output [31:0] io_storeDataQueue_13, // @[:@6.4]
  output [31:0] io_storeDataQueue_14, // @[:@6.4]
  output [31:0] io_storeDataQueue_15, // @[:@6.4]
  input         io_storeDataEnable_0, // @[:@6.4]
  input  [31:0] io_dataFromStorePorts_0, // @[:@6.4]
  input         io_storeAddrEnable_0, // @[:@6.4]
  input  [30:0] io_addressFromStorePorts_0, // @[:@6.4]
  output [30:0] io_storeAddrToMem, // @[:@6.4]
  output [31:0] io_storeDataToMem, // @[:@6.4]
  input         io_storeQIdxOut_ready, // @[:@6.4]
  output        io_storeQIdxOut_valid, // @[:@6.4]
  output [3:0]  io_storeQIdxOut_bits, // @[:@6.4]
  input  [3:0]  io_storeQIdxIn, // @[:@6.4]
  input         io_storeQIdxInValid // @[:@6.4]
);
  reg [3:0] dummyHead; // @[AxiStoreQueue.scala 51:26:@8.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[AxiStoreQueue.scala 53:21:@10.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[AxiStoreQueue.scala 55:24:@28.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[AxiStoreQueue.scala 56:22:@46.4]
  reg [31:0] _RAND_33;
  reg [30:0] addrQ_0; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_34;
  reg [30:0] addrQ_1; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_35;
  reg [30:0] addrQ_2; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_36;
  reg [30:0] addrQ_3; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_37;
  reg [30:0] addrQ_4; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_38;
  reg [30:0] addrQ_5; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_39;
  reg [30:0] addrQ_6; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_40;
  reg [30:0] addrQ_7; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_41;
  reg [30:0] addrQ_8; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_42;
  reg [30:0] addrQ_9; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_43;
  reg [30:0] addrQ_10; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_44;
  reg [30:0] addrQ_11; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_45;
  reg [30:0] addrQ_12; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_46;
  reg [30:0] addrQ_13; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_47;
  reg [30:0] addrQ_14; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_48;
  reg [30:0] addrQ_15; // @[AxiStoreQueue.scala 57:22:@64.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[AxiStoreQueue.scala 58:22:@82.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[AxiStoreQueue.scala 59:26:@100.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[AxiStoreQueue.scala 60:26:@118.4]
  reg [31:0] _RAND_97;
  reg  allocatedEntries_0; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_98;
  reg  allocatedEntries_1; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_99;
  reg  allocatedEntries_2; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_100;
  reg  allocatedEntries_3; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_101;
  reg  allocatedEntries_4; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_102;
  reg  allocatedEntries_5; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_103;
  reg  allocatedEntries_6; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_104;
  reg  allocatedEntries_7; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_105;
  reg  allocatedEntries_8; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_106;
  reg  allocatedEntries_9; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_107;
  reg  allocatedEntries_10; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_108;
  reg  allocatedEntries_11; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_109;
  reg  allocatedEntries_12; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_110;
  reg  allocatedEntries_13; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_111;
  reg  allocatedEntries_14; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_112;
  reg  allocatedEntries_15; // @[AxiStoreQueue.scala 61:33:@136.4]
  reg [31:0] _RAND_113;
  reg  storeCompleted_0; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_114;
  reg  storeCompleted_1; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_115;
  reg  storeCompleted_2; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_116;
  reg  storeCompleted_3; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_117;
  reg  storeCompleted_4; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_118;
  reg  storeCompleted_5; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_119;
  reg  storeCompleted_6; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_120;
  reg  storeCompleted_7; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_121;
  reg  storeCompleted_8; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_122;
  reg  storeCompleted_9; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_123;
  reg  storeCompleted_10; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_124;
  reg  storeCompleted_11; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_125;
  reg  storeCompleted_12; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_126;
  reg  storeCompleted_13; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_127;
  reg  storeCompleted_14; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_128;
  reg  storeCompleted_15; // @[AxiStoreQueue.scala 62:31:@154.4]
  reg [31:0] _RAND_129;
  reg  checkBits_0; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_130;
  reg  checkBits_1; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_131;
  reg  checkBits_2; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_132;
  reg  checkBits_3; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_133;
  reg  checkBits_4; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_134;
  reg  checkBits_5; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_135;
  reg  checkBits_6; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_136;
  reg  checkBits_7; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_137;
  reg  checkBits_8; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_138;
  reg  checkBits_9; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_139;
  reg  checkBits_10; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_140;
  reg  checkBits_11; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_141;
  reg  checkBits_12; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_142;
  reg  checkBits_13; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_143;
  reg  checkBits_14; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_144;
  reg  checkBits_15; // @[AxiStoreQueue.scala 63:26:@172.4]
  reg [31:0] _RAND_145;
  wire [5:0] _GEN_1155; // @[util.scala 14:20:@174.4]
  wire [6:0] _T_1604; // @[util.scala 14:20:@174.4]
  wire [6:0] _T_1605; // @[util.scala 14:20:@175.4]
  wire [5:0] _T_1606; // @[util.scala 14:20:@176.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@177.4]
  wire [4:0] _T_1607; // @[util.scala 14:25:@177.4]
  wire [4:0] _GEN_1156; // @[AxiStoreQueue.scala 72:46:@178.4]
  wire  _T_1608; // @[AxiStoreQueue.scala 72:46:@178.4]
  wire  initBits_0; // @[AxiStoreQueue.scala 72:64:@179.4]
  wire [6:0] _T_1613; // @[util.scala 14:20:@181.4]
  wire [6:0] _T_1614; // @[util.scala 14:20:@182.4]
  wire [5:0] _T_1615; // @[util.scala 14:20:@183.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@184.4]
  wire [4:0] _T_1616; // @[util.scala 14:25:@184.4]
  wire  _T_1617; // @[AxiStoreQueue.scala 72:46:@185.4]
  wire  initBits_1; // @[AxiStoreQueue.scala 72:64:@186.4]
  wire [6:0] _T_1622; // @[util.scala 14:20:@188.4]
  wire [6:0] _T_1623; // @[util.scala 14:20:@189.4]
  wire [5:0] _T_1624; // @[util.scala 14:20:@190.4]
  wire [5:0] _GEN_17; // @[util.scala 14:25:@191.4]
  wire [4:0] _T_1625; // @[util.scala 14:25:@191.4]
  wire  _T_1626; // @[AxiStoreQueue.scala 72:46:@192.4]
  wire  initBits_2; // @[AxiStoreQueue.scala 72:64:@193.4]
  wire [6:0] _T_1631; // @[util.scala 14:20:@195.4]
  wire [6:0] _T_1632; // @[util.scala 14:20:@196.4]
  wire [5:0] _T_1633; // @[util.scala 14:20:@197.4]
  wire [5:0] _GEN_18; // @[util.scala 14:25:@198.4]
  wire [4:0] _T_1634; // @[util.scala 14:25:@198.4]
  wire  _T_1635; // @[AxiStoreQueue.scala 72:46:@199.4]
  wire  initBits_3; // @[AxiStoreQueue.scala 72:64:@200.4]
  wire [6:0] _T_1640; // @[util.scala 14:20:@202.4]
  wire [6:0] _T_1641; // @[util.scala 14:20:@203.4]
  wire [5:0] _T_1642; // @[util.scala 14:20:@204.4]
  wire [5:0] _GEN_19; // @[util.scala 14:25:@205.4]
  wire [4:0] _T_1643; // @[util.scala 14:25:@205.4]
  wire  _T_1644; // @[AxiStoreQueue.scala 72:46:@206.4]
  wire  initBits_4; // @[AxiStoreQueue.scala 72:64:@207.4]
  wire [6:0] _T_1649; // @[util.scala 14:20:@209.4]
  wire [6:0] _T_1650; // @[util.scala 14:20:@210.4]
  wire [5:0] _T_1651; // @[util.scala 14:20:@211.4]
  wire [5:0] _GEN_20; // @[util.scala 14:25:@212.4]
  wire [4:0] _T_1652; // @[util.scala 14:25:@212.4]
  wire  _T_1653; // @[AxiStoreQueue.scala 72:46:@213.4]
  wire  initBits_5; // @[AxiStoreQueue.scala 72:64:@214.4]
  wire [6:0] _T_1658; // @[util.scala 14:20:@216.4]
  wire [6:0] _T_1659; // @[util.scala 14:20:@217.4]
  wire [5:0] _T_1660; // @[util.scala 14:20:@218.4]
  wire [5:0] _GEN_21; // @[util.scala 14:25:@219.4]
  wire [4:0] _T_1661; // @[util.scala 14:25:@219.4]
  wire  _T_1662; // @[AxiStoreQueue.scala 72:46:@220.4]
  wire  initBits_6; // @[AxiStoreQueue.scala 72:64:@221.4]
  wire [6:0] _T_1667; // @[util.scala 14:20:@223.4]
  wire [6:0] _T_1668; // @[util.scala 14:20:@224.4]
  wire [5:0] _T_1669; // @[util.scala 14:20:@225.4]
  wire [5:0] _GEN_22; // @[util.scala 14:25:@226.4]
  wire [4:0] _T_1670; // @[util.scala 14:25:@226.4]
  wire  _T_1671; // @[AxiStoreQueue.scala 72:46:@227.4]
  wire  initBits_7; // @[AxiStoreQueue.scala 72:64:@228.4]
  wire [6:0] _T_1676; // @[util.scala 14:20:@230.4]
  wire [6:0] _T_1677; // @[util.scala 14:20:@231.4]
  wire [5:0] _T_1678; // @[util.scala 14:20:@232.4]
  wire [5:0] _GEN_23; // @[util.scala 14:25:@233.4]
  wire [4:0] _T_1679; // @[util.scala 14:25:@233.4]
  wire  _T_1680; // @[AxiStoreQueue.scala 72:46:@234.4]
  wire  initBits_8; // @[AxiStoreQueue.scala 72:64:@235.4]
  wire [6:0] _T_1685; // @[util.scala 14:20:@237.4]
  wire [6:0] _T_1686; // @[util.scala 14:20:@238.4]
  wire [5:0] _T_1687; // @[util.scala 14:20:@239.4]
  wire [5:0] _GEN_24; // @[util.scala 14:25:@240.4]
  wire [4:0] _T_1688; // @[util.scala 14:25:@240.4]
  wire  _T_1689; // @[AxiStoreQueue.scala 72:46:@241.4]
  wire  initBits_9; // @[AxiStoreQueue.scala 72:64:@242.4]
  wire [6:0] _T_1694; // @[util.scala 14:20:@244.4]
  wire [6:0] _T_1695; // @[util.scala 14:20:@245.4]
  wire [5:0] _T_1696; // @[util.scala 14:20:@246.4]
  wire [5:0] _GEN_25; // @[util.scala 14:25:@247.4]
  wire [4:0] _T_1697; // @[util.scala 14:25:@247.4]
  wire  _T_1698; // @[AxiStoreQueue.scala 72:46:@248.4]
  wire  initBits_10; // @[AxiStoreQueue.scala 72:64:@249.4]
  wire [6:0] _T_1703; // @[util.scala 14:20:@251.4]
  wire [6:0] _T_1704; // @[util.scala 14:20:@252.4]
  wire [5:0] _T_1705; // @[util.scala 14:20:@253.4]
  wire [5:0] _GEN_26; // @[util.scala 14:25:@254.4]
  wire [4:0] _T_1706; // @[util.scala 14:25:@254.4]
  wire  _T_1707; // @[AxiStoreQueue.scala 72:46:@255.4]
  wire  initBits_11; // @[AxiStoreQueue.scala 72:64:@256.4]
  wire [6:0] _T_1712; // @[util.scala 14:20:@258.4]
  wire [6:0] _T_1713; // @[util.scala 14:20:@259.4]
  wire [5:0] _T_1714; // @[util.scala 14:20:@260.4]
  wire [5:0] _GEN_27; // @[util.scala 14:25:@261.4]
  wire [4:0] _T_1715; // @[util.scala 14:25:@261.4]
  wire  _T_1716; // @[AxiStoreQueue.scala 72:46:@262.4]
  wire  initBits_12; // @[AxiStoreQueue.scala 72:64:@263.4]
  wire [6:0] _T_1721; // @[util.scala 14:20:@265.4]
  wire [6:0] _T_1722; // @[util.scala 14:20:@266.4]
  wire [5:0] _T_1723; // @[util.scala 14:20:@267.4]
  wire [5:0] _GEN_28; // @[util.scala 14:25:@268.4]
  wire [4:0] _T_1724; // @[util.scala 14:25:@268.4]
  wire  _T_1725; // @[AxiStoreQueue.scala 72:46:@269.4]
  wire  initBits_13; // @[AxiStoreQueue.scala 72:64:@270.4]
  wire [6:0] _T_1730; // @[util.scala 14:20:@272.4]
  wire [6:0] _T_1731; // @[util.scala 14:20:@273.4]
  wire [5:0] _T_1732; // @[util.scala 14:20:@274.4]
  wire [5:0] _GEN_29; // @[util.scala 14:25:@275.4]
  wire [4:0] _T_1733; // @[util.scala 14:25:@275.4]
  wire  _T_1734; // @[AxiStoreQueue.scala 72:46:@276.4]
  wire  initBits_14; // @[AxiStoreQueue.scala 72:64:@277.4]
  wire [6:0] _T_1739; // @[util.scala 14:20:@279.4]
  wire [6:0] _T_1740; // @[util.scala 14:20:@280.4]
  wire [5:0] _T_1741; // @[util.scala 14:20:@281.4]
  wire [5:0] _GEN_30; // @[util.scala 14:25:@282.4]
  wire [4:0] _T_1742; // @[util.scala 14:25:@282.4]
  wire  _T_1743; // @[AxiStoreQueue.scala 72:46:@283.4]
  wire  initBits_15; // @[AxiStoreQueue.scala 72:64:@284.4]
  wire  _T_1766; // @[AxiStoreQueue.scala 74:78:@302.4]
  wire  _T_1767; // @[AxiStoreQueue.scala 74:78:@303.4]
  wire  _T_1768; // @[AxiStoreQueue.scala 74:78:@304.4]
  wire  _T_1769; // @[AxiStoreQueue.scala 74:78:@305.4]
  wire  _T_1770; // @[AxiStoreQueue.scala 74:78:@306.4]
  wire  _T_1771; // @[AxiStoreQueue.scala 74:78:@307.4]
  wire  _T_1772; // @[AxiStoreQueue.scala 74:78:@308.4]
  wire  _T_1773; // @[AxiStoreQueue.scala 74:78:@309.4]
  wire  _T_1774; // @[AxiStoreQueue.scala 74:78:@310.4]
  wire  _T_1775; // @[AxiStoreQueue.scala 74:78:@311.4]
  wire  _T_1776; // @[AxiStoreQueue.scala 74:78:@312.4]
  wire  _T_1777; // @[AxiStoreQueue.scala 74:78:@313.4]
  wire  _T_1778; // @[AxiStoreQueue.scala 74:78:@314.4]
  wire  _T_1779; // @[AxiStoreQueue.scala 74:78:@315.4]
  wire  _T_1780; // @[AxiStoreQueue.scala 74:78:@316.4]
  wire  _T_1781; // @[AxiStoreQueue.scala 74:78:@317.4]
  wire [3:0] _T_1812; // @[:@357.6]
  wire [3:0] _GEN_1; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_2; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_3; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_4; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_5; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_6; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_7; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_8; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_9; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_10; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_11; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_12; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_13; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_14; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_15; // @[AxiStoreQueue.scala 78:20:@358.6]
  wire [3:0] _GEN_32; // @[AxiStoreQueue.scala 77:25:@351.4]
  wire  _GEN_33; // @[AxiStoreQueue.scala 77:25:@351.4]
  wire [3:0] _T_1830; // @[:@373.6]
  wire [3:0] _GEN_35; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_36; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_37; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_38; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_39; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_40; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_41; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_42; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_43; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_44; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_45; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_46; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_47; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_48; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_49; // @[AxiStoreQueue.scala 78:20:@374.6]
  wire [3:0] _GEN_66; // @[AxiStoreQueue.scala 77:25:@367.4]
  wire  _GEN_67; // @[AxiStoreQueue.scala 77:25:@367.4]
  wire [3:0] _T_1848; // @[:@389.6]
  wire [3:0] _GEN_69; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_70; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_71; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_72; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_73; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_74; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_75; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_76; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_77; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_78; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_79; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_80; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_81; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_82; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_83; // @[AxiStoreQueue.scala 78:20:@390.6]
  wire [3:0] _GEN_100; // @[AxiStoreQueue.scala 77:25:@383.4]
  wire  _GEN_101; // @[AxiStoreQueue.scala 77:25:@383.4]
  wire [3:0] _T_1866; // @[:@405.6]
  wire [3:0] _GEN_103; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_104; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_105; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_106; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_107; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_108; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_109; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_110; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_111; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_112; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_113; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_114; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_115; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_116; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_117; // @[AxiStoreQueue.scala 78:20:@406.6]
  wire [3:0] _GEN_134; // @[AxiStoreQueue.scala 77:25:@399.4]
  wire  _GEN_135; // @[AxiStoreQueue.scala 77:25:@399.4]
  wire [3:0] _T_1884; // @[:@421.6]
  wire [3:0] _GEN_137; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_138; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_139; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_140; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_141; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_142; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_143; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_144; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_145; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_146; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_147; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_148; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_149; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_150; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_151; // @[AxiStoreQueue.scala 78:20:@422.6]
  wire [3:0] _GEN_168; // @[AxiStoreQueue.scala 77:25:@415.4]
  wire  _GEN_169; // @[AxiStoreQueue.scala 77:25:@415.4]
  wire [3:0] _T_1902; // @[:@437.6]
  wire [3:0] _GEN_171; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_172; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_173; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_174; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_175; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_176; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_177; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_178; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_179; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_180; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_181; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_182; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_183; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_184; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_185; // @[AxiStoreQueue.scala 78:20:@438.6]
  wire [3:0] _GEN_202; // @[AxiStoreQueue.scala 77:25:@431.4]
  wire  _GEN_203; // @[AxiStoreQueue.scala 77:25:@431.4]
  wire [3:0] _T_1920; // @[:@453.6]
  wire [3:0] _GEN_205; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_206; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_207; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_208; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_209; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_210; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_211; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_212; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_213; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_214; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_215; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_216; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_217; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_218; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_219; // @[AxiStoreQueue.scala 78:20:@454.6]
  wire [3:0] _GEN_236; // @[AxiStoreQueue.scala 77:25:@447.4]
  wire  _GEN_237; // @[AxiStoreQueue.scala 77:25:@447.4]
  wire [3:0] _T_1938; // @[:@469.6]
  wire [3:0] _GEN_239; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_240; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_241; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_242; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_243; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_244; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_245; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_246; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_247; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_248; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_249; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_250; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_251; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_252; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_253; // @[AxiStoreQueue.scala 78:20:@470.6]
  wire [3:0] _GEN_270; // @[AxiStoreQueue.scala 77:25:@463.4]
  wire  _GEN_271; // @[AxiStoreQueue.scala 77:25:@463.4]
  wire [3:0] _T_1956; // @[:@485.6]
  wire [3:0] _GEN_273; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_274; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_275; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_276; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_277; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_278; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_279; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_280; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_281; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_282; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_283; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_284; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_285; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_286; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_287; // @[AxiStoreQueue.scala 78:20:@486.6]
  wire [3:0] _GEN_304; // @[AxiStoreQueue.scala 77:25:@479.4]
  wire  _GEN_305; // @[AxiStoreQueue.scala 77:25:@479.4]
  wire [3:0] _T_1974; // @[:@501.6]
  wire [3:0] _GEN_307; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_308; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_309; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_310; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_311; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_312; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_313; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_314; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_315; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_316; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_317; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_318; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_319; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_320; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_321; // @[AxiStoreQueue.scala 78:20:@502.6]
  wire [3:0] _GEN_338; // @[AxiStoreQueue.scala 77:25:@495.4]
  wire  _GEN_339; // @[AxiStoreQueue.scala 77:25:@495.4]
  wire [3:0] _T_1992; // @[:@517.6]
  wire [3:0] _GEN_341; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_342; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_343; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_344; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_345; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_346; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_347; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_348; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_349; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_350; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_351; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_352; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_353; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_354; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_355; // @[AxiStoreQueue.scala 78:20:@518.6]
  wire [3:0] _GEN_372; // @[AxiStoreQueue.scala 77:25:@511.4]
  wire  _GEN_373; // @[AxiStoreQueue.scala 77:25:@511.4]
  wire [3:0] _T_2010; // @[:@533.6]
  wire [3:0] _GEN_375; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_376; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_377; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_378; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_379; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_380; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_381; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_382; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_383; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_384; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_385; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_386; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_387; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_388; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_389; // @[AxiStoreQueue.scala 78:20:@534.6]
  wire [3:0] _GEN_406; // @[AxiStoreQueue.scala 77:25:@527.4]
  wire  _GEN_407; // @[AxiStoreQueue.scala 77:25:@527.4]
  wire [3:0] _T_2028; // @[:@549.6]
  wire [3:0] _GEN_409; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_410; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_411; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_412; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_413; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_414; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_415; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_416; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_417; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_418; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_419; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_420; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_421; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_422; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_423; // @[AxiStoreQueue.scala 78:20:@550.6]
  wire [3:0] _GEN_440; // @[AxiStoreQueue.scala 77:25:@543.4]
  wire  _GEN_441; // @[AxiStoreQueue.scala 77:25:@543.4]
  wire [3:0] _T_2046; // @[:@565.6]
  wire [3:0] _GEN_443; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_444; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_445; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_446; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_447; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_448; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_449; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_450; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_451; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_452; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_453; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_454; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_455; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_456; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_457; // @[AxiStoreQueue.scala 78:20:@566.6]
  wire [3:0] _GEN_474; // @[AxiStoreQueue.scala 77:25:@559.4]
  wire  _GEN_475; // @[AxiStoreQueue.scala 77:25:@559.4]
  wire [3:0] _T_2064; // @[:@581.6]
  wire [3:0] _GEN_477; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_478; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_479; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_480; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_481; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_482; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_483; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_484; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_485; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_486; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_487; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_488; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_489; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_490; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_491; // @[AxiStoreQueue.scala 78:20:@582.6]
  wire [3:0] _GEN_508; // @[AxiStoreQueue.scala 77:25:@575.4]
  wire  _GEN_509; // @[AxiStoreQueue.scala 77:25:@575.4]
  wire [3:0] _T_2082; // @[:@597.6]
  wire [3:0] _GEN_511; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_512; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_513; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_514; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_515; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_516; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_517; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_518; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_519; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_520; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_521; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_522; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_523; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_524; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_525; // @[AxiStoreQueue.scala 78:20:@598.6]
  wire [3:0] _GEN_542; // @[AxiStoreQueue.scala 77:25:@591.4]
  wire  _GEN_543; // @[AxiStoreQueue.scala 77:25:@591.4]
  reg [3:0] previousLoadHead; // @[AxiStoreQueue.scala 94:33:@607.4]
  reg [31:0] _RAND_146;
  wire [4:0] _T_2104; // @[util.scala 10:8:@616.6]
  wire [4:0] _GEN_31; // @[util.scala 10:14:@617.6]
  wire [4:0] _T_2105; // @[util.scala 10:14:@617.6]
  wire [4:0] _GEN_1220; // @[AxiStoreQueue.scala 98:56:@618.6]
  wire  _T_2106; // @[AxiStoreQueue.scala 98:56:@618.6]
  wire  _T_2107; // @[AxiStoreQueue.scala 97:50:@619.6]
  wire  _T_2109; // @[AxiStoreQueue.scala 97:35:@620.6]
  wire  _T_2111; // @[AxiStoreQueue.scala 102:35:@628.8]
  wire  _T_2112; // @[AxiStoreQueue.scala 102:87:@629.8]
  wire  _T_2113; // @[AxiStoreQueue.scala 102:61:@630.8]
  wire  _T_2115; // @[AxiStoreQueue.scala 104:35:@635.10]
  wire  _T_2116; // @[AxiStoreQueue.scala 105:23:@636.10]
  wire  _T_2117; // @[AxiStoreQueue.scala 105:75:@637.10]
  wire  _T_2118; // @[AxiStoreQueue.scala 105:49:@638.10]
  wire  _T_2120; // @[AxiStoreQueue.scala 105:9:@639.10]
  wire  _T_2121; // @[AxiStoreQueue.scala 104:49:@640.10]
  wire  _GEN_560; // @[AxiStoreQueue.scala 105:96:@641.10]
  wire  _GEN_561; // @[AxiStoreQueue.scala 102:102:@631.8]
  wire  _GEN_562; // @[AxiStoreQueue.scala 100:26:@624.6]
  wire  _GEN_563; // @[AxiStoreQueue.scala 96:35:@609.4]
  wire [4:0] _T_2134; // @[util.scala 10:8:@652.6]
  wire [4:0] _GEN_34; // @[util.scala 10:14:@653.6]
  wire [4:0] _T_2135; // @[util.scala 10:14:@653.6]
  wire  _T_2136; // @[AxiStoreQueue.scala 98:56:@654.6]
  wire  _T_2137; // @[AxiStoreQueue.scala 97:50:@655.6]
  wire  _T_2139; // @[AxiStoreQueue.scala 97:35:@656.6]
  wire  _T_2141; // @[AxiStoreQueue.scala 102:35:@664.8]
  wire  _T_2142; // @[AxiStoreQueue.scala 102:87:@665.8]
  wire  _T_2143; // @[AxiStoreQueue.scala 102:61:@666.8]
  wire  _T_2146; // @[AxiStoreQueue.scala 105:23:@672.10]
  wire  _T_2147; // @[AxiStoreQueue.scala 105:75:@673.10]
  wire  _T_2148; // @[AxiStoreQueue.scala 105:49:@674.10]
  wire  _T_2150; // @[AxiStoreQueue.scala 105:9:@675.10]
  wire  _T_2151; // @[AxiStoreQueue.scala 104:49:@676.10]
  wire  _GEN_580; // @[AxiStoreQueue.scala 105:96:@677.10]
  wire  _GEN_581; // @[AxiStoreQueue.scala 102:102:@667.8]
  wire  _GEN_582; // @[AxiStoreQueue.scala 100:26:@660.6]
  wire  _GEN_583; // @[AxiStoreQueue.scala 96:35:@645.4]
  wire [4:0] _T_2164; // @[util.scala 10:8:@688.6]
  wire [4:0] _GEN_50; // @[util.scala 10:14:@689.6]
  wire [4:0] _T_2165; // @[util.scala 10:14:@689.6]
  wire  _T_2166; // @[AxiStoreQueue.scala 98:56:@690.6]
  wire  _T_2167; // @[AxiStoreQueue.scala 97:50:@691.6]
  wire  _T_2169; // @[AxiStoreQueue.scala 97:35:@692.6]
  wire  _T_2171; // @[AxiStoreQueue.scala 102:35:@700.8]
  wire  _T_2172; // @[AxiStoreQueue.scala 102:87:@701.8]
  wire  _T_2173; // @[AxiStoreQueue.scala 102:61:@702.8]
  wire  _T_2176; // @[AxiStoreQueue.scala 105:23:@708.10]
  wire  _T_2177; // @[AxiStoreQueue.scala 105:75:@709.10]
  wire  _T_2178; // @[AxiStoreQueue.scala 105:49:@710.10]
  wire  _T_2180; // @[AxiStoreQueue.scala 105:9:@711.10]
  wire  _T_2181; // @[AxiStoreQueue.scala 104:49:@712.10]
  wire  _GEN_600; // @[AxiStoreQueue.scala 105:96:@713.10]
  wire  _GEN_601; // @[AxiStoreQueue.scala 102:102:@703.8]
  wire  _GEN_602; // @[AxiStoreQueue.scala 100:26:@696.6]
  wire  _GEN_603; // @[AxiStoreQueue.scala 96:35:@681.4]
  wire [4:0] _T_2194; // @[util.scala 10:8:@724.6]
  wire [4:0] _GEN_51; // @[util.scala 10:14:@725.6]
  wire [4:0] _T_2195; // @[util.scala 10:14:@725.6]
  wire  _T_2196; // @[AxiStoreQueue.scala 98:56:@726.6]
  wire  _T_2197; // @[AxiStoreQueue.scala 97:50:@727.6]
  wire  _T_2199; // @[AxiStoreQueue.scala 97:35:@728.6]
  wire  _T_2201; // @[AxiStoreQueue.scala 102:35:@736.8]
  wire  _T_2202; // @[AxiStoreQueue.scala 102:87:@737.8]
  wire  _T_2203; // @[AxiStoreQueue.scala 102:61:@738.8]
  wire  _T_2206; // @[AxiStoreQueue.scala 105:23:@744.10]
  wire  _T_2207; // @[AxiStoreQueue.scala 105:75:@745.10]
  wire  _T_2208; // @[AxiStoreQueue.scala 105:49:@746.10]
  wire  _T_2210; // @[AxiStoreQueue.scala 105:9:@747.10]
  wire  _T_2211; // @[AxiStoreQueue.scala 104:49:@748.10]
  wire  _GEN_620; // @[AxiStoreQueue.scala 105:96:@749.10]
  wire  _GEN_621; // @[AxiStoreQueue.scala 102:102:@739.8]
  wire  _GEN_622; // @[AxiStoreQueue.scala 100:26:@732.6]
  wire  _GEN_623; // @[AxiStoreQueue.scala 96:35:@717.4]
  wire [4:0] _T_2224; // @[util.scala 10:8:@760.6]
  wire [4:0] _GEN_52; // @[util.scala 10:14:@761.6]
  wire [4:0] _T_2225; // @[util.scala 10:14:@761.6]
  wire  _T_2226; // @[AxiStoreQueue.scala 98:56:@762.6]
  wire  _T_2227; // @[AxiStoreQueue.scala 97:50:@763.6]
  wire  _T_2229; // @[AxiStoreQueue.scala 97:35:@764.6]
  wire  _T_2231; // @[AxiStoreQueue.scala 102:35:@772.8]
  wire  _T_2232; // @[AxiStoreQueue.scala 102:87:@773.8]
  wire  _T_2233; // @[AxiStoreQueue.scala 102:61:@774.8]
  wire  _T_2236; // @[AxiStoreQueue.scala 105:23:@780.10]
  wire  _T_2237; // @[AxiStoreQueue.scala 105:75:@781.10]
  wire  _T_2238; // @[AxiStoreQueue.scala 105:49:@782.10]
  wire  _T_2240; // @[AxiStoreQueue.scala 105:9:@783.10]
  wire  _T_2241; // @[AxiStoreQueue.scala 104:49:@784.10]
  wire  _GEN_640; // @[AxiStoreQueue.scala 105:96:@785.10]
  wire  _GEN_641; // @[AxiStoreQueue.scala 102:102:@775.8]
  wire  _GEN_642; // @[AxiStoreQueue.scala 100:26:@768.6]
  wire  _GEN_643; // @[AxiStoreQueue.scala 96:35:@753.4]
  wire [4:0] _T_2254; // @[util.scala 10:8:@796.6]
  wire [4:0] _GEN_53; // @[util.scala 10:14:@797.6]
  wire [4:0] _T_2255; // @[util.scala 10:14:@797.6]
  wire  _T_2256; // @[AxiStoreQueue.scala 98:56:@798.6]
  wire  _T_2257; // @[AxiStoreQueue.scala 97:50:@799.6]
  wire  _T_2259; // @[AxiStoreQueue.scala 97:35:@800.6]
  wire  _T_2261; // @[AxiStoreQueue.scala 102:35:@808.8]
  wire  _T_2262; // @[AxiStoreQueue.scala 102:87:@809.8]
  wire  _T_2263; // @[AxiStoreQueue.scala 102:61:@810.8]
  wire  _T_2266; // @[AxiStoreQueue.scala 105:23:@816.10]
  wire  _T_2267; // @[AxiStoreQueue.scala 105:75:@817.10]
  wire  _T_2268; // @[AxiStoreQueue.scala 105:49:@818.10]
  wire  _T_2270; // @[AxiStoreQueue.scala 105:9:@819.10]
  wire  _T_2271; // @[AxiStoreQueue.scala 104:49:@820.10]
  wire  _GEN_660; // @[AxiStoreQueue.scala 105:96:@821.10]
  wire  _GEN_661; // @[AxiStoreQueue.scala 102:102:@811.8]
  wire  _GEN_662; // @[AxiStoreQueue.scala 100:26:@804.6]
  wire  _GEN_663; // @[AxiStoreQueue.scala 96:35:@789.4]
  wire [4:0] _T_2284; // @[util.scala 10:8:@832.6]
  wire [4:0] _GEN_54; // @[util.scala 10:14:@833.6]
  wire [4:0] _T_2285; // @[util.scala 10:14:@833.6]
  wire  _T_2286; // @[AxiStoreQueue.scala 98:56:@834.6]
  wire  _T_2287; // @[AxiStoreQueue.scala 97:50:@835.6]
  wire  _T_2289; // @[AxiStoreQueue.scala 97:35:@836.6]
  wire  _T_2291; // @[AxiStoreQueue.scala 102:35:@844.8]
  wire  _T_2292; // @[AxiStoreQueue.scala 102:87:@845.8]
  wire  _T_2293; // @[AxiStoreQueue.scala 102:61:@846.8]
  wire  _T_2296; // @[AxiStoreQueue.scala 105:23:@852.10]
  wire  _T_2297; // @[AxiStoreQueue.scala 105:75:@853.10]
  wire  _T_2298; // @[AxiStoreQueue.scala 105:49:@854.10]
  wire  _T_2300; // @[AxiStoreQueue.scala 105:9:@855.10]
  wire  _T_2301; // @[AxiStoreQueue.scala 104:49:@856.10]
  wire  _GEN_680; // @[AxiStoreQueue.scala 105:96:@857.10]
  wire  _GEN_681; // @[AxiStoreQueue.scala 102:102:@847.8]
  wire  _GEN_682; // @[AxiStoreQueue.scala 100:26:@840.6]
  wire  _GEN_683; // @[AxiStoreQueue.scala 96:35:@825.4]
  wire [4:0] _T_2314; // @[util.scala 10:8:@868.6]
  wire [4:0] _GEN_55; // @[util.scala 10:14:@869.6]
  wire [4:0] _T_2315; // @[util.scala 10:14:@869.6]
  wire  _T_2316; // @[AxiStoreQueue.scala 98:56:@870.6]
  wire  _T_2317; // @[AxiStoreQueue.scala 97:50:@871.6]
  wire  _T_2319; // @[AxiStoreQueue.scala 97:35:@872.6]
  wire  _T_2321; // @[AxiStoreQueue.scala 102:35:@880.8]
  wire  _T_2322; // @[AxiStoreQueue.scala 102:87:@881.8]
  wire  _T_2323; // @[AxiStoreQueue.scala 102:61:@882.8]
  wire  _T_2326; // @[AxiStoreQueue.scala 105:23:@888.10]
  wire  _T_2327; // @[AxiStoreQueue.scala 105:75:@889.10]
  wire  _T_2328; // @[AxiStoreQueue.scala 105:49:@890.10]
  wire  _T_2330; // @[AxiStoreQueue.scala 105:9:@891.10]
  wire  _T_2331; // @[AxiStoreQueue.scala 104:49:@892.10]
  wire  _GEN_700; // @[AxiStoreQueue.scala 105:96:@893.10]
  wire  _GEN_701; // @[AxiStoreQueue.scala 102:102:@883.8]
  wire  _GEN_702; // @[AxiStoreQueue.scala 100:26:@876.6]
  wire  _GEN_703; // @[AxiStoreQueue.scala 96:35:@861.4]
  wire [4:0] _T_2344; // @[util.scala 10:8:@904.6]
  wire [4:0] _GEN_56; // @[util.scala 10:14:@905.6]
  wire [4:0] _T_2345; // @[util.scala 10:14:@905.6]
  wire  _T_2346; // @[AxiStoreQueue.scala 98:56:@906.6]
  wire  _T_2347; // @[AxiStoreQueue.scala 97:50:@907.6]
  wire  _T_2349; // @[AxiStoreQueue.scala 97:35:@908.6]
  wire  _T_2351; // @[AxiStoreQueue.scala 102:35:@916.8]
  wire  _T_2352; // @[AxiStoreQueue.scala 102:87:@917.8]
  wire  _T_2353; // @[AxiStoreQueue.scala 102:61:@918.8]
  wire  _T_2356; // @[AxiStoreQueue.scala 105:23:@924.10]
  wire  _T_2357; // @[AxiStoreQueue.scala 105:75:@925.10]
  wire  _T_2358; // @[AxiStoreQueue.scala 105:49:@926.10]
  wire  _T_2360; // @[AxiStoreQueue.scala 105:9:@927.10]
  wire  _T_2361; // @[AxiStoreQueue.scala 104:49:@928.10]
  wire  _GEN_720; // @[AxiStoreQueue.scala 105:96:@929.10]
  wire  _GEN_721; // @[AxiStoreQueue.scala 102:102:@919.8]
  wire  _GEN_722; // @[AxiStoreQueue.scala 100:26:@912.6]
  wire  _GEN_723; // @[AxiStoreQueue.scala 96:35:@897.4]
  wire [4:0] _T_2374; // @[util.scala 10:8:@940.6]
  wire [4:0] _GEN_57; // @[util.scala 10:14:@941.6]
  wire [4:0] _T_2375; // @[util.scala 10:14:@941.6]
  wire  _T_2376; // @[AxiStoreQueue.scala 98:56:@942.6]
  wire  _T_2377; // @[AxiStoreQueue.scala 97:50:@943.6]
  wire  _T_2379; // @[AxiStoreQueue.scala 97:35:@944.6]
  wire  _T_2381; // @[AxiStoreQueue.scala 102:35:@952.8]
  wire  _T_2382; // @[AxiStoreQueue.scala 102:87:@953.8]
  wire  _T_2383; // @[AxiStoreQueue.scala 102:61:@954.8]
  wire  _T_2386; // @[AxiStoreQueue.scala 105:23:@960.10]
  wire  _T_2387; // @[AxiStoreQueue.scala 105:75:@961.10]
  wire  _T_2388; // @[AxiStoreQueue.scala 105:49:@962.10]
  wire  _T_2390; // @[AxiStoreQueue.scala 105:9:@963.10]
  wire  _T_2391; // @[AxiStoreQueue.scala 104:49:@964.10]
  wire  _GEN_740; // @[AxiStoreQueue.scala 105:96:@965.10]
  wire  _GEN_741; // @[AxiStoreQueue.scala 102:102:@955.8]
  wire  _GEN_742; // @[AxiStoreQueue.scala 100:26:@948.6]
  wire  _GEN_743; // @[AxiStoreQueue.scala 96:35:@933.4]
  wire [4:0] _T_2404; // @[util.scala 10:8:@976.6]
  wire [4:0] _GEN_58; // @[util.scala 10:14:@977.6]
  wire [4:0] _T_2405; // @[util.scala 10:14:@977.6]
  wire  _T_2406; // @[AxiStoreQueue.scala 98:56:@978.6]
  wire  _T_2407; // @[AxiStoreQueue.scala 97:50:@979.6]
  wire  _T_2409; // @[AxiStoreQueue.scala 97:35:@980.6]
  wire  _T_2411; // @[AxiStoreQueue.scala 102:35:@988.8]
  wire  _T_2412; // @[AxiStoreQueue.scala 102:87:@989.8]
  wire  _T_2413; // @[AxiStoreQueue.scala 102:61:@990.8]
  wire  _T_2416; // @[AxiStoreQueue.scala 105:23:@996.10]
  wire  _T_2417; // @[AxiStoreQueue.scala 105:75:@997.10]
  wire  _T_2418; // @[AxiStoreQueue.scala 105:49:@998.10]
  wire  _T_2420; // @[AxiStoreQueue.scala 105:9:@999.10]
  wire  _T_2421; // @[AxiStoreQueue.scala 104:49:@1000.10]
  wire  _GEN_760; // @[AxiStoreQueue.scala 105:96:@1001.10]
  wire  _GEN_761; // @[AxiStoreQueue.scala 102:102:@991.8]
  wire  _GEN_762; // @[AxiStoreQueue.scala 100:26:@984.6]
  wire  _GEN_763; // @[AxiStoreQueue.scala 96:35:@969.4]
  wire [4:0] _T_2434; // @[util.scala 10:8:@1012.6]
  wire [4:0] _GEN_59; // @[util.scala 10:14:@1013.6]
  wire [4:0] _T_2435; // @[util.scala 10:14:@1013.6]
  wire  _T_2436; // @[AxiStoreQueue.scala 98:56:@1014.6]
  wire  _T_2437; // @[AxiStoreQueue.scala 97:50:@1015.6]
  wire  _T_2439; // @[AxiStoreQueue.scala 97:35:@1016.6]
  wire  _T_2441; // @[AxiStoreQueue.scala 102:35:@1024.8]
  wire  _T_2442; // @[AxiStoreQueue.scala 102:87:@1025.8]
  wire  _T_2443; // @[AxiStoreQueue.scala 102:61:@1026.8]
  wire  _T_2446; // @[AxiStoreQueue.scala 105:23:@1032.10]
  wire  _T_2447; // @[AxiStoreQueue.scala 105:75:@1033.10]
  wire  _T_2448; // @[AxiStoreQueue.scala 105:49:@1034.10]
  wire  _T_2450; // @[AxiStoreQueue.scala 105:9:@1035.10]
  wire  _T_2451; // @[AxiStoreQueue.scala 104:49:@1036.10]
  wire  _GEN_780; // @[AxiStoreQueue.scala 105:96:@1037.10]
  wire  _GEN_781; // @[AxiStoreQueue.scala 102:102:@1027.8]
  wire  _GEN_782; // @[AxiStoreQueue.scala 100:26:@1020.6]
  wire  _GEN_783; // @[AxiStoreQueue.scala 96:35:@1005.4]
  wire [4:0] _T_2464; // @[util.scala 10:8:@1048.6]
  wire [4:0] _GEN_60; // @[util.scala 10:14:@1049.6]
  wire [4:0] _T_2465; // @[util.scala 10:14:@1049.6]
  wire  _T_2466; // @[AxiStoreQueue.scala 98:56:@1050.6]
  wire  _T_2467; // @[AxiStoreQueue.scala 97:50:@1051.6]
  wire  _T_2469; // @[AxiStoreQueue.scala 97:35:@1052.6]
  wire  _T_2471; // @[AxiStoreQueue.scala 102:35:@1060.8]
  wire  _T_2472; // @[AxiStoreQueue.scala 102:87:@1061.8]
  wire  _T_2473; // @[AxiStoreQueue.scala 102:61:@1062.8]
  wire  _T_2476; // @[AxiStoreQueue.scala 105:23:@1068.10]
  wire  _T_2477; // @[AxiStoreQueue.scala 105:75:@1069.10]
  wire  _T_2478; // @[AxiStoreQueue.scala 105:49:@1070.10]
  wire  _T_2480; // @[AxiStoreQueue.scala 105:9:@1071.10]
  wire  _T_2481; // @[AxiStoreQueue.scala 104:49:@1072.10]
  wire  _GEN_800; // @[AxiStoreQueue.scala 105:96:@1073.10]
  wire  _GEN_801; // @[AxiStoreQueue.scala 102:102:@1063.8]
  wire  _GEN_802; // @[AxiStoreQueue.scala 100:26:@1056.6]
  wire  _GEN_803; // @[AxiStoreQueue.scala 96:35:@1041.4]
  wire [4:0] _T_2494; // @[util.scala 10:8:@1084.6]
  wire [4:0] _GEN_61; // @[util.scala 10:14:@1085.6]
  wire [4:0] _T_2495; // @[util.scala 10:14:@1085.6]
  wire  _T_2496; // @[AxiStoreQueue.scala 98:56:@1086.6]
  wire  _T_2497; // @[AxiStoreQueue.scala 97:50:@1087.6]
  wire  _T_2499; // @[AxiStoreQueue.scala 97:35:@1088.6]
  wire  _T_2501; // @[AxiStoreQueue.scala 102:35:@1096.8]
  wire  _T_2502; // @[AxiStoreQueue.scala 102:87:@1097.8]
  wire  _T_2503; // @[AxiStoreQueue.scala 102:61:@1098.8]
  wire  _T_2506; // @[AxiStoreQueue.scala 105:23:@1104.10]
  wire  _T_2507; // @[AxiStoreQueue.scala 105:75:@1105.10]
  wire  _T_2508; // @[AxiStoreQueue.scala 105:49:@1106.10]
  wire  _T_2510; // @[AxiStoreQueue.scala 105:9:@1107.10]
  wire  _T_2511; // @[AxiStoreQueue.scala 104:49:@1108.10]
  wire  _GEN_820; // @[AxiStoreQueue.scala 105:96:@1109.10]
  wire  _GEN_821; // @[AxiStoreQueue.scala 102:102:@1099.8]
  wire  _GEN_822; // @[AxiStoreQueue.scala 100:26:@1092.6]
  wire  _GEN_823; // @[AxiStoreQueue.scala 96:35:@1077.4]
  wire [4:0] _T_2524; // @[util.scala 10:8:@1120.6]
  wire [4:0] _GEN_62; // @[util.scala 10:14:@1121.6]
  wire [4:0] _T_2525; // @[util.scala 10:14:@1121.6]
  wire  _T_2526; // @[AxiStoreQueue.scala 98:56:@1122.6]
  wire  _T_2527; // @[AxiStoreQueue.scala 97:50:@1123.6]
  wire  _T_2529; // @[AxiStoreQueue.scala 97:35:@1124.6]
  wire  _T_2531; // @[AxiStoreQueue.scala 102:35:@1132.8]
  wire  _T_2532; // @[AxiStoreQueue.scala 102:87:@1133.8]
  wire  _T_2533; // @[AxiStoreQueue.scala 102:61:@1134.8]
  wire  _T_2536; // @[AxiStoreQueue.scala 105:23:@1140.10]
  wire  _T_2537; // @[AxiStoreQueue.scala 105:75:@1141.10]
  wire  _T_2538; // @[AxiStoreQueue.scala 105:49:@1142.10]
  wire  _T_2540; // @[AxiStoreQueue.scala 105:9:@1143.10]
  wire  _T_2541; // @[AxiStoreQueue.scala 104:49:@1144.10]
  wire  _GEN_840; // @[AxiStoreQueue.scala 105:96:@1145.10]
  wire  _GEN_841; // @[AxiStoreQueue.scala 102:102:@1135.8]
  wire  _GEN_842; // @[AxiStoreQueue.scala 100:26:@1128.6]
  wire  _GEN_843; // @[AxiStoreQueue.scala 96:35:@1113.4]
  wire [4:0] _T_2554; // @[util.scala 10:8:@1156.6]
  wire [4:0] _GEN_63; // @[util.scala 10:14:@1157.6]
  wire [4:0] _T_2555; // @[util.scala 10:14:@1157.6]
  wire  _T_2556; // @[AxiStoreQueue.scala 98:56:@1158.6]
  wire  _T_2557; // @[AxiStoreQueue.scala 97:50:@1159.6]
  wire  _T_2559; // @[AxiStoreQueue.scala 97:35:@1160.6]
  wire  _T_2561; // @[AxiStoreQueue.scala 102:35:@1168.8]
  wire  _T_2562; // @[AxiStoreQueue.scala 102:87:@1169.8]
  wire  _T_2563; // @[AxiStoreQueue.scala 102:61:@1170.8]
  wire  _T_2566; // @[AxiStoreQueue.scala 105:23:@1176.10]
  wire  _T_2567; // @[AxiStoreQueue.scala 105:75:@1177.10]
  wire  _T_2568; // @[AxiStoreQueue.scala 105:49:@1178.10]
  wire  _T_2570; // @[AxiStoreQueue.scala 105:9:@1179.10]
  wire  _T_2571; // @[AxiStoreQueue.scala 104:49:@1180.10]
  wire  _GEN_860; // @[AxiStoreQueue.scala 105:96:@1181.10]
  wire  _GEN_861; // @[AxiStoreQueue.scala 102:102:@1171.8]
  wire  _GEN_862; // @[AxiStoreQueue.scala 100:26:@1164.6]
  wire  _GEN_863; // @[AxiStoreQueue.scala 96:35:@1149.4]
  wire  _T_2573; // @[AxiStoreQueue.scala 121:103:@1185.4]
  wire  _T_2575; // @[AxiStoreQueue.scala 122:17:@1186.4]
  wire  _T_2577; // @[AxiStoreQueue.scala 122:35:@1187.4]
  wire  _T_2578; // @[AxiStoreQueue.scala 122:26:@1188.4]
  wire  _T_2580; // @[AxiStoreQueue.scala 122:50:@1189.4]
  wire  _T_2582; // @[AxiStoreQueue.scala 122:81:@1190.4]
  wire  _T_2584; // @[AxiStoreQueue.scala 122:99:@1191.4]
  wire  _T_2585; // @[AxiStoreQueue.scala 122:90:@1192.4]
  wire  _T_2587; // @[AxiStoreQueue.scala 122:67:@1193.4]
  wire  _T_2588; // @[AxiStoreQueue.scala 122:64:@1194.4]
  wire  validEntriesInLoadQ_0; // @[AxiStoreQueue.scala 121:90:@1195.4]
  wire  _T_2592; // @[AxiStoreQueue.scala 122:17:@1197.4]
  wire  _T_2594; // @[AxiStoreQueue.scala 122:35:@1198.4]
  wire  _T_2595; // @[AxiStoreQueue.scala 122:26:@1199.4]
  wire  _T_2599; // @[AxiStoreQueue.scala 122:81:@1201.4]
  wire  _T_2601; // @[AxiStoreQueue.scala 122:99:@1202.4]
  wire  _T_2602; // @[AxiStoreQueue.scala 122:90:@1203.4]
  wire  _T_2604; // @[AxiStoreQueue.scala 122:67:@1204.4]
  wire  _T_2605; // @[AxiStoreQueue.scala 122:64:@1205.4]
  wire  validEntriesInLoadQ_1; // @[AxiStoreQueue.scala 121:90:@1206.4]
  wire  _T_2609; // @[AxiStoreQueue.scala 122:17:@1208.4]
  wire  _T_2611; // @[AxiStoreQueue.scala 122:35:@1209.4]
  wire  _T_2612; // @[AxiStoreQueue.scala 122:26:@1210.4]
  wire  _T_2616; // @[AxiStoreQueue.scala 122:81:@1212.4]
  wire  _T_2618; // @[AxiStoreQueue.scala 122:99:@1213.4]
  wire  _T_2619; // @[AxiStoreQueue.scala 122:90:@1214.4]
  wire  _T_2621; // @[AxiStoreQueue.scala 122:67:@1215.4]
  wire  _T_2622; // @[AxiStoreQueue.scala 122:64:@1216.4]
  wire  validEntriesInLoadQ_2; // @[AxiStoreQueue.scala 121:90:@1217.4]
  wire  _T_2626; // @[AxiStoreQueue.scala 122:17:@1219.4]
  wire  _T_2628; // @[AxiStoreQueue.scala 122:35:@1220.4]
  wire  _T_2629; // @[AxiStoreQueue.scala 122:26:@1221.4]
  wire  _T_2633; // @[AxiStoreQueue.scala 122:81:@1223.4]
  wire  _T_2635; // @[AxiStoreQueue.scala 122:99:@1224.4]
  wire  _T_2636; // @[AxiStoreQueue.scala 122:90:@1225.4]
  wire  _T_2638; // @[AxiStoreQueue.scala 122:67:@1226.4]
  wire  _T_2639; // @[AxiStoreQueue.scala 122:64:@1227.4]
  wire  validEntriesInLoadQ_3; // @[AxiStoreQueue.scala 121:90:@1228.4]
  wire  _T_2643; // @[AxiStoreQueue.scala 122:17:@1230.4]
  wire  _T_2645; // @[AxiStoreQueue.scala 122:35:@1231.4]
  wire  _T_2646; // @[AxiStoreQueue.scala 122:26:@1232.4]
  wire  _T_2650; // @[AxiStoreQueue.scala 122:81:@1234.4]
  wire  _T_2652; // @[AxiStoreQueue.scala 122:99:@1235.4]
  wire  _T_2653; // @[AxiStoreQueue.scala 122:90:@1236.4]
  wire  _T_2655; // @[AxiStoreQueue.scala 122:67:@1237.4]
  wire  _T_2656; // @[AxiStoreQueue.scala 122:64:@1238.4]
  wire  validEntriesInLoadQ_4; // @[AxiStoreQueue.scala 121:90:@1239.4]
  wire  _T_2660; // @[AxiStoreQueue.scala 122:17:@1241.4]
  wire  _T_2662; // @[AxiStoreQueue.scala 122:35:@1242.4]
  wire  _T_2663; // @[AxiStoreQueue.scala 122:26:@1243.4]
  wire  _T_2667; // @[AxiStoreQueue.scala 122:81:@1245.4]
  wire  _T_2669; // @[AxiStoreQueue.scala 122:99:@1246.4]
  wire  _T_2670; // @[AxiStoreQueue.scala 122:90:@1247.4]
  wire  _T_2672; // @[AxiStoreQueue.scala 122:67:@1248.4]
  wire  _T_2673; // @[AxiStoreQueue.scala 122:64:@1249.4]
  wire  validEntriesInLoadQ_5; // @[AxiStoreQueue.scala 121:90:@1250.4]
  wire  _T_2677; // @[AxiStoreQueue.scala 122:17:@1252.4]
  wire  _T_2679; // @[AxiStoreQueue.scala 122:35:@1253.4]
  wire  _T_2680; // @[AxiStoreQueue.scala 122:26:@1254.4]
  wire  _T_2684; // @[AxiStoreQueue.scala 122:81:@1256.4]
  wire  _T_2686; // @[AxiStoreQueue.scala 122:99:@1257.4]
  wire  _T_2687; // @[AxiStoreQueue.scala 122:90:@1258.4]
  wire  _T_2689; // @[AxiStoreQueue.scala 122:67:@1259.4]
  wire  _T_2690; // @[AxiStoreQueue.scala 122:64:@1260.4]
  wire  validEntriesInLoadQ_6; // @[AxiStoreQueue.scala 121:90:@1261.4]
  wire  _T_2694; // @[AxiStoreQueue.scala 122:17:@1263.4]
  wire  _T_2696; // @[AxiStoreQueue.scala 122:35:@1264.4]
  wire  _T_2697; // @[AxiStoreQueue.scala 122:26:@1265.4]
  wire  _T_2701; // @[AxiStoreQueue.scala 122:81:@1267.4]
  wire  _T_2703; // @[AxiStoreQueue.scala 122:99:@1268.4]
  wire  _T_2704; // @[AxiStoreQueue.scala 122:90:@1269.4]
  wire  _T_2706; // @[AxiStoreQueue.scala 122:67:@1270.4]
  wire  _T_2707; // @[AxiStoreQueue.scala 122:64:@1271.4]
  wire  validEntriesInLoadQ_7; // @[AxiStoreQueue.scala 121:90:@1272.4]
  wire  _T_2711; // @[AxiStoreQueue.scala 122:17:@1274.4]
  wire  _T_2713; // @[AxiStoreQueue.scala 122:35:@1275.4]
  wire  _T_2714; // @[AxiStoreQueue.scala 122:26:@1276.4]
  wire  _T_2718; // @[AxiStoreQueue.scala 122:81:@1278.4]
  wire  _T_2720; // @[AxiStoreQueue.scala 122:99:@1279.4]
  wire  _T_2721; // @[AxiStoreQueue.scala 122:90:@1280.4]
  wire  _T_2723; // @[AxiStoreQueue.scala 122:67:@1281.4]
  wire  _T_2724; // @[AxiStoreQueue.scala 122:64:@1282.4]
  wire  validEntriesInLoadQ_8; // @[AxiStoreQueue.scala 121:90:@1283.4]
  wire  _T_2728; // @[AxiStoreQueue.scala 122:17:@1285.4]
  wire  _T_2730; // @[AxiStoreQueue.scala 122:35:@1286.4]
  wire  _T_2731; // @[AxiStoreQueue.scala 122:26:@1287.4]
  wire  _T_2735; // @[AxiStoreQueue.scala 122:81:@1289.4]
  wire  _T_2737; // @[AxiStoreQueue.scala 122:99:@1290.4]
  wire  _T_2738; // @[AxiStoreQueue.scala 122:90:@1291.4]
  wire  _T_2740; // @[AxiStoreQueue.scala 122:67:@1292.4]
  wire  _T_2741; // @[AxiStoreQueue.scala 122:64:@1293.4]
  wire  validEntriesInLoadQ_9; // @[AxiStoreQueue.scala 121:90:@1294.4]
  wire  _T_2745; // @[AxiStoreQueue.scala 122:17:@1296.4]
  wire  _T_2747; // @[AxiStoreQueue.scala 122:35:@1297.4]
  wire  _T_2748; // @[AxiStoreQueue.scala 122:26:@1298.4]
  wire  _T_2752; // @[AxiStoreQueue.scala 122:81:@1300.4]
  wire  _T_2754; // @[AxiStoreQueue.scala 122:99:@1301.4]
  wire  _T_2755; // @[AxiStoreQueue.scala 122:90:@1302.4]
  wire  _T_2757; // @[AxiStoreQueue.scala 122:67:@1303.4]
  wire  _T_2758; // @[AxiStoreQueue.scala 122:64:@1304.4]
  wire  validEntriesInLoadQ_10; // @[AxiStoreQueue.scala 121:90:@1305.4]
  wire  _T_2762; // @[AxiStoreQueue.scala 122:17:@1307.4]
  wire  _T_2764; // @[AxiStoreQueue.scala 122:35:@1308.4]
  wire  _T_2765; // @[AxiStoreQueue.scala 122:26:@1309.4]
  wire  _T_2769; // @[AxiStoreQueue.scala 122:81:@1311.4]
  wire  _T_2771; // @[AxiStoreQueue.scala 122:99:@1312.4]
  wire  _T_2772; // @[AxiStoreQueue.scala 122:90:@1313.4]
  wire  _T_2774; // @[AxiStoreQueue.scala 122:67:@1314.4]
  wire  _T_2775; // @[AxiStoreQueue.scala 122:64:@1315.4]
  wire  validEntriesInLoadQ_11; // @[AxiStoreQueue.scala 121:90:@1316.4]
  wire  _T_2779; // @[AxiStoreQueue.scala 122:17:@1318.4]
  wire  _T_2781; // @[AxiStoreQueue.scala 122:35:@1319.4]
  wire  _T_2782; // @[AxiStoreQueue.scala 122:26:@1320.4]
  wire  _T_2786; // @[AxiStoreQueue.scala 122:81:@1322.4]
  wire  _T_2788; // @[AxiStoreQueue.scala 122:99:@1323.4]
  wire  _T_2789; // @[AxiStoreQueue.scala 122:90:@1324.4]
  wire  _T_2791; // @[AxiStoreQueue.scala 122:67:@1325.4]
  wire  _T_2792; // @[AxiStoreQueue.scala 122:64:@1326.4]
  wire  validEntriesInLoadQ_12; // @[AxiStoreQueue.scala 121:90:@1327.4]
  wire  _T_2796; // @[AxiStoreQueue.scala 122:17:@1329.4]
  wire  _T_2798; // @[AxiStoreQueue.scala 122:35:@1330.4]
  wire  _T_2799; // @[AxiStoreQueue.scala 122:26:@1331.4]
  wire  _T_2803; // @[AxiStoreQueue.scala 122:81:@1333.4]
  wire  _T_2805; // @[AxiStoreQueue.scala 122:99:@1334.4]
  wire  _T_2806; // @[AxiStoreQueue.scala 122:90:@1335.4]
  wire  _T_2808; // @[AxiStoreQueue.scala 122:67:@1336.4]
  wire  _T_2809; // @[AxiStoreQueue.scala 122:64:@1337.4]
  wire  validEntriesInLoadQ_13; // @[AxiStoreQueue.scala 121:90:@1338.4]
  wire  _T_2813; // @[AxiStoreQueue.scala 122:17:@1340.4]
  wire  _T_2815; // @[AxiStoreQueue.scala 122:35:@1341.4]
  wire  _T_2816; // @[AxiStoreQueue.scala 122:26:@1342.4]
  wire  _T_2820; // @[AxiStoreQueue.scala 122:81:@1344.4]
  wire  _T_2822; // @[AxiStoreQueue.scala 122:99:@1345.4]
  wire  _T_2823; // @[AxiStoreQueue.scala 122:90:@1346.4]
  wire  _T_2825; // @[AxiStoreQueue.scala 122:67:@1347.4]
  wire  _T_2826; // @[AxiStoreQueue.scala 122:64:@1348.4]
  wire  validEntriesInLoadQ_14; // @[AxiStoreQueue.scala 121:90:@1349.4]
  wire  validEntriesInLoadQ_15; // @[AxiStoreQueue.scala 121:90:@1360.4]
  wire [3:0] _GEN_865; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_866; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_867; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_868; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_869; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_870; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_871; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_872; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_873; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_874; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_875; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_876; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_877; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_878; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire [3:0] _GEN_879; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire  _T_2869; // @[AxiStoreQueue.scala 128:96:@1378.4]
  wire  loadsToCheck_0; // @[AxiStoreQueue.scala 128:83:@1386.4]
  wire  _T_2899; // @[AxiStoreQueue.scala 129:35:@1389.4]
  wire  _T_2900; // @[AxiStoreQueue.scala 129:26:@1390.4]
  wire  _T_2905; // @[AxiStoreQueue.scala 129:79:@1391.4]
  wire  _T_2908; // @[AxiStoreQueue.scala 129:87:@1393.4]
  wire  _T_2910; // @[AxiStoreQueue.scala 129:58:@1394.4]
  wire  loadsToCheck_1; // @[AxiStoreQueue.scala 128:83:@1395.4]
  wire  _T_2922; // @[AxiStoreQueue.scala 129:35:@1398.4]
  wire  _T_2923; // @[AxiStoreQueue.scala 129:26:@1399.4]
  wire  _T_2928; // @[AxiStoreQueue.scala 129:79:@1400.4]
  wire  _T_2931; // @[AxiStoreQueue.scala 129:87:@1402.4]
  wire  _T_2933; // @[AxiStoreQueue.scala 129:58:@1403.4]
  wire  loadsToCheck_2; // @[AxiStoreQueue.scala 128:83:@1404.4]
  wire  _T_2945; // @[AxiStoreQueue.scala 129:35:@1407.4]
  wire  _T_2946; // @[AxiStoreQueue.scala 129:26:@1408.4]
  wire  _T_2951; // @[AxiStoreQueue.scala 129:79:@1409.4]
  wire  _T_2954; // @[AxiStoreQueue.scala 129:87:@1411.4]
  wire  _T_2956; // @[AxiStoreQueue.scala 129:58:@1412.4]
  wire  loadsToCheck_3; // @[AxiStoreQueue.scala 128:83:@1413.4]
  wire  _T_2968; // @[AxiStoreQueue.scala 129:35:@1416.4]
  wire  _T_2969; // @[AxiStoreQueue.scala 129:26:@1417.4]
  wire  _T_2974; // @[AxiStoreQueue.scala 129:79:@1418.4]
  wire  _T_2977; // @[AxiStoreQueue.scala 129:87:@1420.4]
  wire  _T_2979; // @[AxiStoreQueue.scala 129:58:@1421.4]
  wire  loadsToCheck_4; // @[AxiStoreQueue.scala 128:83:@1422.4]
  wire  _T_2991; // @[AxiStoreQueue.scala 129:35:@1425.4]
  wire  _T_2992; // @[AxiStoreQueue.scala 129:26:@1426.4]
  wire  _T_2997; // @[AxiStoreQueue.scala 129:79:@1427.4]
  wire  _T_3000; // @[AxiStoreQueue.scala 129:87:@1429.4]
  wire  _T_3002; // @[AxiStoreQueue.scala 129:58:@1430.4]
  wire  loadsToCheck_5; // @[AxiStoreQueue.scala 128:83:@1431.4]
  wire  _T_3014; // @[AxiStoreQueue.scala 129:35:@1434.4]
  wire  _T_3015; // @[AxiStoreQueue.scala 129:26:@1435.4]
  wire  _T_3020; // @[AxiStoreQueue.scala 129:79:@1436.4]
  wire  _T_3023; // @[AxiStoreQueue.scala 129:87:@1438.4]
  wire  _T_3025; // @[AxiStoreQueue.scala 129:58:@1439.4]
  wire  loadsToCheck_6; // @[AxiStoreQueue.scala 128:83:@1440.4]
  wire  _T_3037; // @[AxiStoreQueue.scala 129:35:@1443.4]
  wire  _T_3038; // @[AxiStoreQueue.scala 129:26:@1444.4]
  wire  _T_3043; // @[AxiStoreQueue.scala 129:79:@1445.4]
  wire  _T_3046; // @[AxiStoreQueue.scala 129:87:@1447.4]
  wire  _T_3048; // @[AxiStoreQueue.scala 129:58:@1448.4]
  wire  loadsToCheck_7; // @[AxiStoreQueue.scala 128:83:@1449.4]
  wire  _T_3060; // @[AxiStoreQueue.scala 129:35:@1452.4]
  wire  _T_3061; // @[AxiStoreQueue.scala 129:26:@1453.4]
  wire  _T_3066; // @[AxiStoreQueue.scala 129:79:@1454.4]
  wire  _T_3069; // @[AxiStoreQueue.scala 129:87:@1456.4]
  wire  _T_3071; // @[AxiStoreQueue.scala 129:58:@1457.4]
  wire  loadsToCheck_8; // @[AxiStoreQueue.scala 128:83:@1458.4]
  wire  _T_3083; // @[AxiStoreQueue.scala 129:35:@1461.4]
  wire  _T_3084; // @[AxiStoreQueue.scala 129:26:@1462.4]
  wire  _T_3089; // @[AxiStoreQueue.scala 129:79:@1463.4]
  wire  _T_3092; // @[AxiStoreQueue.scala 129:87:@1465.4]
  wire  _T_3094; // @[AxiStoreQueue.scala 129:58:@1466.4]
  wire  loadsToCheck_9; // @[AxiStoreQueue.scala 128:83:@1467.4]
  wire  _T_3106; // @[AxiStoreQueue.scala 129:35:@1470.4]
  wire  _T_3107; // @[AxiStoreQueue.scala 129:26:@1471.4]
  wire  _T_3112; // @[AxiStoreQueue.scala 129:79:@1472.4]
  wire  _T_3115; // @[AxiStoreQueue.scala 129:87:@1474.4]
  wire  _T_3117; // @[AxiStoreQueue.scala 129:58:@1475.4]
  wire  loadsToCheck_10; // @[AxiStoreQueue.scala 128:83:@1476.4]
  wire  _T_3129; // @[AxiStoreQueue.scala 129:35:@1479.4]
  wire  _T_3130; // @[AxiStoreQueue.scala 129:26:@1480.4]
  wire  _T_3135; // @[AxiStoreQueue.scala 129:79:@1481.4]
  wire  _T_3138; // @[AxiStoreQueue.scala 129:87:@1483.4]
  wire  _T_3140; // @[AxiStoreQueue.scala 129:58:@1484.4]
  wire  loadsToCheck_11; // @[AxiStoreQueue.scala 128:83:@1485.4]
  wire  _T_3152; // @[AxiStoreQueue.scala 129:35:@1488.4]
  wire  _T_3153; // @[AxiStoreQueue.scala 129:26:@1489.4]
  wire  _T_3158; // @[AxiStoreQueue.scala 129:79:@1490.4]
  wire  _T_3161; // @[AxiStoreQueue.scala 129:87:@1492.4]
  wire  _T_3163; // @[AxiStoreQueue.scala 129:58:@1493.4]
  wire  loadsToCheck_12; // @[AxiStoreQueue.scala 128:83:@1494.4]
  wire  _T_3175; // @[AxiStoreQueue.scala 129:35:@1497.4]
  wire  _T_3176; // @[AxiStoreQueue.scala 129:26:@1498.4]
  wire  _T_3181; // @[AxiStoreQueue.scala 129:79:@1499.4]
  wire  _T_3184; // @[AxiStoreQueue.scala 129:87:@1501.4]
  wire  _T_3186; // @[AxiStoreQueue.scala 129:58:@1502.4]
  wire  loadsToCheck_13; // @[AxiStoreQueue.scala 128:83:@1503.4]
  wire  _T_3198; // @[AxiStoreQueue.scala 129:35:@1506.4]
  wire  _T_3199; // @[AxiStoreQueue.scala 129:26:@1507.4]
  wire  _T_3204; // @[AxiStoreQueue.scala 129:79:@1508.4]
  wire  _T_3207; // @[AxiStoreQueue.scala 129:87:@1510.4]
  wire  _T_3209; // @[AxiStoreQueue.scala 129:58:@1511.4]
  wire  loadsToCheck_14; // @[AxiStoreQueue.scala 128:83:@1512.4]
  wire  _T_3221; // @[AxiStoreQueue.scala 129:35:@1515.4]
  wire  loadsToCheck_15; // @[AxiStoreQueue.scala 128:83:@1521.4]
  wire  _T_3255; // @[AxiStoreQueue.scala 135:16:@1539.4]
  wire  _GEN_881; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_882; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_883; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_884; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_885; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_886; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_887; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_888; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_889; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_890; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_891; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_892; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_893; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_894; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _GEN_895; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  entriesToCheck_0; // @[AxiStoreQueue.scala 135:24:@1540.4]
  wire  _T_3260; // @[AxiStoreQueue.scala 135:16:@1541.4]
  wire  entriesToCheck_1; // @[AxiStoreQueue.scala 135:24:@1542.4]
  wire  _T_3265; // @[AxiStoreQueue.scala 135:16:@1543.4]
  wire  entriesToCheck_2; // @[AxiStoreQueue.scala 135:24:@1544.4]
  wire  _T_3270; // @[AxiStoreQueue.scala 135:16:@1545.4]
  wire  entriesToCheck_3; // @[AxiStoreQueue.scala 135:24:@1546.4]
  wire  _T_3275; // @[AxiStoreQueue.scala 135:16:@1547.4]
  wire  entriesToCheck_4; // @[AxiStoreQueue.scala 135:24:@1548.4]
  wire  _T_3280; // @[AxiStoreQueue.scala 135:16:@1549.4]
  wire  entriesToCheck_5; // @[AxiStoreQueue.scala 135:24:@1550.4]
  wire  _T_3285; // @[AxiStoreQueue.scala 135:16:@1551.4]
  wire  entriesToCheck_6; // @[AxiStoreQueue.scala 135:24:@1552.4]
  wire  _T_3290; // @[AxiStoreQueue.scala 135:16:@1553.4]
  wire  entriesToCheck_7; // @[AxiStoreQueue.scala 135:24:@1554.4]
  wire  _T_3295; // @[AxiStoreQueue.scala 135:16:@1555.4]
  wire  entriesToCheck_8; // @[AxiStoreQueue.scala 135:24:@1556.4]
  wire  _T_3300; // @[AxiStoreQueue.scala 135:16:@1557.4]
  wire  entriesToCheck_9; // @[AxiStoreQueue.scala 135:24:@1558.4]
  wire  _T_3305; // @[AxiStoreQueue.scala 135:16:@1559.4]
  wire  entriesToCheck_10; // @[AxiStoreQueue.scala 135:24:@1560.4]
  wire  _T_3310; // @[AxiStoreQueue.scala 135:16:@1561.4]
  wire  entriesToCheck_11; // @[AxiStoreQueue.scala 135:24:@1562.4]
  wire  _T_3315; // @[AxiStoreQueue.scala 135:16:@1563.4]
  wire  entriesToCheck_12; // @[AxiStoreQueue.scala 135:24:@1564.4]
  wire  _T_3320; // @[AxiStoreQueue.scala 135:16:@1565.4]
  wire  entriesToCheck_13; // @[AxiStoreQueue.scala 135:24:@1566.4]
  wire  _T_3325; // @[AxiStoreQueue.scala 135:16:@1567.4]
  wire  entriesToCheck_14; // @[AxiStoreQueue.scala 135:24:@1568.4]
  wire  _T_3330; // @[AxiStoreQueue.scala 135:16:@1569.4]
  wire  entriesToCheck_15; // @[AxiStoreQueue.scala 135:24:@1570.4]
  wire  _T_3378; // @[AxiStoreQueue.scala 142:34:@1589.4]
  wire  _T_3379; // @[AxiStoreQueue.scala 142:64:@1590.4]
  wire [30:0] _GEN_897; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_898; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_899; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_900; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_901; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_902; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_903; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_904; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_905; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_906; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_907; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_908; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_909; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_910; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire [30:0] _GEN_911; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire  _T_3383; // @[AxiStoreQueue.scala 143:56:@1591.4]
  wire  _T_3384; // @[AxiStoreQueue.scala 143:36:@1592.4]
  wire  noConflicts_0; // @[AxiStoreQueue.scala 142:95:@1593.4]
  wire  _T_3387; // @[AxiStoreQueue.scala 142:34:@1595.4]
  wire  _T_3388; // @[AxiStoreQueue.scala 142:64:@1596.4]
  wire  _T_3392; // @[AxiStoreQueue.scala 143:56:@1597.4]
  wire  _T_3393; // @[AxiStoreQueue.scala 143:36:@1598.4]
  wire  noConflicts_1; // @[AxiStoreQueue.scala 142:95:@1599.4]
  wire  _T_3396; // @[AxiStoreQueue.scala 142:34:@1601.4]
  wire  _T_3397; // @[AxiStoreQueue.scala 142:64:@1602.4]
  wire  _T_3401; // @[AxiStoreQueue.scala 143:56:@1603.4]
  wire  _T_3402; // @[AxiStoreQueue.scala 143:36:@1604.4]
  wire  noConflicts_2; // @[AxiStoreQueue.scala 142:95:@1605.4]
  wire  _T_3405; // @[AxiStoreQueue.scala 142:34:@1607.4]
  wire  _T_3406; // @[AxiStoreQueue.scala 142:64:@1608.4]
  wire  _T_3410; // @[AxiStoreQueue.scala 143:56:@1609.4]
  wire  _T_3411; // @[AxiStoreQueue.scala 143:36:@1610.4]
  wire  noConflicts_3; // @[AxiStoreQueue.scala 142:95:@1611.4]
  wire  _T_3414; // @[AxiStoreQueue.scala 142:34:@1613.4]
  wire  _T_3415; // @[AxiStoreQueue.scala 142:64:@1614.4]
  wire  _T_3419; // @[AxiStoreQueue.scala 143:56:@1615.4]
  wire  _T_3420; // @[AxiStoreQueue.scala 143:36:@1616.4]
  wire  noConflicts_4; // @[AxiStoreQueue.scala 142:95:@1617.4]
  wire  _T_3423; // @[AxiStoreQueue.scala 142:34:@1619.4]
  wire  _T_3424; // @[AxiStoreQueue.scala 142:64:@1620.4]
  wire  _T_3428; // @[AxiStoreQueue.scala 143:56:@1621.4]
  wire  _T_3429; // @[AxiStoreQueue.scala 143:36:@1622.4]
  wire  noConflicts_5; // @[AxiStoreQueue.scala 142:95:@1623.4]
  wire  _T_3432; // @[AxiStoreQueue.scala 142:34:@1625.4]
  wire  _T_3433; // @[AxiStoreQueue.scala 142:64:@1626.4]
  wire  _T_3437; // @[AxiStoreQueue.scala 143:56:@1627.4]
  wire  _T_3438; // @[AxiStoreQueue.scala 143:36:@1628.4]
  wire  noConflicts_6; // @[AxiStoreQueue.scala 142:95:@1629.4]
  wire  _T_3441; // @[AxiStoreQueue.scala 142:34:@1631.4]
  wire  _T_3442; // @[AxiStoreQueue.scala 142:64:@1632.4]
  wire  _T_3446; // @[AxiStoreQueue.scala 143:56:@1633.4]
  wire  _T_3447; // @[AxiStoreQueue.scala 143:36:@1634.4]
  wire  noConflicts_7; // @[AxiStoreQueue.scala 142:95:@1635.4]
  wire  _T_3450; // @[AxiStoreQueue.scala 142:34:@1637.4]
  wire  _T_3451; // @[AxiStoreQueue.scala 142:64:@1638.4]
  wire  _T_3455; // @[AxiStoreQueue.scala 143:56:@1639.4]
  wire  _T_3456; // @[AxiStoreQueue.scala 143:36:@1640.4]
  wire  noConflicts_8; // @[AxiStoreQueue.scala 142:95:@1641.4]
  wire  _T_3459; // @[AxiStoreQueue.scala 142:34:@1643.4]
  wire  _T_3460; // @[AxiStoreQueue.scala 142:64:@1644.4]
  wire  _T_3464; // @[AxiStoreQueue.scala 143:56:@1645.4]
  wire  _T_3465; // @[AxiStoreQueue.scala 143:36:@1646.4]
  wire  noConflicts_9; // @[AxiStoreQueue.scala 142:95:@1647.4]
  wire  _T_3468; // @[AxiStoreQueue.scala 142:34:@1649.4]
  wire  _T_3469; // @[AxiStoreQueue.scala 142:64:@1650.4]
  wire  _T_3473; // @[AxiStoreQueue.scala 143:56:@1651.4]
  wire  _T_3474; // @[AxiStoreQueue.scala 143:36:@1652.4]
  wire  noConflicts_10; // @[AxiStoreQueue.scala 142:95:@1653.4]
  wire  _T_3477; // @[AxiStoreQueue.scala 142:34:@1655.4]
  wire  _T_3478; // @[AxiStoreQueue.scala 142:64:@1656.4]
  wire  _T_3482; // @[AxiStoreQueue.scala 143:56:@1657.4]
  wire  _T_3483; // @[AxiStoreQueue.scala 143:36:@1658.4]
  wire  noConflicts_11; // @[AxiStoreQueue.scala 142:95:@1659.4]
  wire  _T_3486; // @[AxiStoreQueue.scala 142:34:@1661.4]
  wire  _T_3487; // @[AxiStoreQueue.scala 142:64:@1662.4]
  wire  _T_3491; // @[AxiStoreQueue.scala 143:56:@1663.4]
  wire  _T_3492; // @[AxiStoreQueue.scala 143:36:@1664.4]
  wire  noConflicts_12; // @[AxiStoreQueue.scala 142:95:@1665.4]
  wire  _T_3495; // @[AxiStoreQueue.scala 142:34:@1667.4]
  wire  _T_3496; // @[AxiStoreQueue.scala 142:64:@1668.4]
  wire  _T_3500; // @[AxiStoreQueue.scala 143:56:@1669.4]
  wire  _T_3501; // @[AxiStoreQueue.scala 143:36:@1670.4]
  wire  noConflicts_13; // @[AxiStoreQueue.scala 142:95:@1671.4]
  wire  _T_3504; // @[AxiStoreQueue.scala 142:34:@1673.4]
  wire  _T_3505; // @[AxiStoreQueue.scala 142:64:@1674.4]
  wire  _T_3509; // @[AxiStoreQueue.scala 143:56:@1675.4]
  wire  _T_3510; // @[AxiStoreQueue.scala 143:36:@1676.4]
  wire  noConflicts_14; // @[AxiStoreQueue.scala 142:95:@1677.4]
  wire  _T_3513; // @[AxiStoreQueue.scala 142:34:@1679.4]
  wire  _T_3514; // @[AxiStoreQueue.scala 142:64:@1680.4]
  wire  _T_3518; // @[AxiStoreQueue.scala 143:56:@1681.4]
  wire  _T_3519; // @[AxiStoreQueue.scala 143:36:@1682.4]
  wire  noConflicts_15; // @[AxiStoreQueue.scala 142:95:@1683.4]
  wire  _GEN_913; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_914; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_915; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_916; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_917; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_918; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_919; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_920; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_921; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_922; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_923; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_924; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_925; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_926; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_927; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_929; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_930; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_931; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_932; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_933; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_934; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_935; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_936; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_937; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_938; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_939; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_940; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_941; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_942; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_943; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _T_3527; // @[AxiStoreQueue.scala 156:49:@1685.4]
  wire  _GEN_945; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_946; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_947; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_948; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_949; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_950; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_951; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_952; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_953; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_954; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_955; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_956; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_957; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_958; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _GEN_959; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _T_3532; // @[AxiStoreQueue.scala 156:76:@1686.4]
  wire  _T_3533; // @[AxiStoreQueue.scala 156:73:@1687.4]
  wire  _T_3536; // @[AxiStoreQueue.scala 156:124:@1689.4]
  wire  _T_3537; // @[AxiStoreQueue.scala 156:124:@1690.4]
  wire  _T_3538; // @[AxiStoreQueue.scala 156:124:@1691.4]
  wire  _T_3539; // @[AxiStoreQueue.scala 156:124:@1692.4]
  wire  _T_3540; // @[AxiStoreQueue.scala 156:124:@1693.4]
  wire  _T_3541; // @[AxiStoreQueue.scala 156:124:@1694.4]
  wire  _T_3542; // @[AxiStoreQueue.scala 156:124:@1695.4]
  wire  _T_3543; // @[AxiStoreQueue.scala 156:124:@1696.4]
  wire  _T_3544; // @[AxiStoreQueue.scala 156:124:@1697.4]
  wire  _T_3545; // @[AxiStoreQueue.scala 156:124:@1698.4]
  wire  _T_3546; // @[AxiStoreQueue.scala 156:124:@1699.4]
  wire  _T_3547; // @[AxiStoreQueue.scala 156:124:@1700.4]
  wire  _T_3548; // @[AxiStoreQueue.scala 156:124:@1701.4]
  wire  _T_3549; // @[AxiStoreQueue.scala 156:124:@1702.4]
  wire  _T_3550; // @[AxiStoreQueue.scala 156:124:@1703.4]
  wire  storeRequest; // @[AxiStoreQueue.scala 156:103:@1704.4]
  wire  _T_3553; // @[AxiStoreQueue.scala 168:54:@1710.6]
  wire  _T_3554; // @[AxiStoreQueue.scala 168:36:@1711.6]
  wire  _GEN_960; // @[AxiStoreQueue.scala 168:75:@1712.6]
  wire  _GEN_961; // @[AxiStoreQueue.scala 166:35:@1706.4]
  wire  _T_3558; // @[AxiStoreQueue.scala 168:54:@1719.6]
  wire  _T_3559; // @[AxiStoreQueue.scala 168:36:@1720.6]
  wire  _GEN_962; // @[AxiStoreQueue.scala 168:75:@1721.6]
  wire  _GEN_963; // @[AxiStoreQueue.scala 166:35:@1715.4]
  wire  _T_3563; // @[AxiStoreQueue.scala 168:54:@1728.6]
  wire  _T_3564; // @[AxiStoreQueue.scala 168:36:@1729.6]
  wire  _GEN_964; // @[AxiStoreQueue.scala 168:75:@1730.6]
  wire  _GEN_965; // @[AxiStoreQueue.scala 166:35:@1724.4]
  wire  _T_3568; // @[AxiStoreQueue.scala 168:54:@1737.6]
  wire  _T_3569; // @[AxiStoreQueue.scala 168:36:@1738.6]
  wire  _GEN_966; // @[AxiStoreQueue.scala 168:75:@1739.6]
  wire  _GEN_967; // @[AxiStoreQueue.scala 166:35:@1733.4]
  wire  _T_3573; // @[AxiStoreQueue.scala 168:54:@1746.6]
  wire  _T_3574; // @[AxiStoreQueue.scala 168:36:@1747.6]
  wire  _GEN_968; // @[AxiStoreQueue.scala 168:75:@1748.6]
  wire  _GEN_969; // @[AxiStoreQueue.scala 166:35:@1742.4]
  wire  _T_3578; // @[AxiStoreQueue.scala 168:54:@1755.6]
  wire  _T_3579; // @[AxiStoreQueue.scala 168:36:@1756.6]
  wire  _GEN_970; // @[AxiStoreQueue.scala 168:75:@1757.6]
  wire  _GEN_971; // @[AxiStoreQueue.scala 166:35:@1751.4]
  wire  _T_3583; // @[AxiStoreQueue.scala 168:54:@1764.6]
  wire  _T_3584; // @[AxiStoreQueue.scala 168:36:@1765.6]
  wire  _GEN_972; // @[AxiStoreQueue.scala 168:75:@1766.6]
  wire  _GEN_973; // @[AxiStoreQueue.scala 166:35:@1760.4]
  wire  _T_3588; // @[AxiStoreQueue.scala 168:54:@1773.6]
  wire  _T_3589; // @[AxiStoreQueue.scala 168:36:@1774.6]
  wire  _GEN_974; // @[AxiStoreQueue.scala 168:75:@1775.6]
  wire  _GEN_975; // @[AxiStoreQueue.scala 166:35:@1769.4]
  wire  _T_3593; // @[AxiStoreQueue.scala 168:54:@1782.6]
  wire  _T_3594; // @[AxiStoreQueue.scala 168:36:@1783.6]
  wire  _GEN_976; // @[AxiStoreQueue.scala 168:75:@1784.6]
  wire  _GEN_977; // @[AxiStoreQueue.scala 166:35:@1778.4]
  wire  _T_3598; // @[AxiStoreQueue.scala 168:54:@1791.6]
  wire  _T_3599; // @[AxiStoreQueue.scala 168:36:@1792.6]
  wire  _GEN_978; // @[AxiStoreQueue.scala 168:75:@1793.6]
  wire  _GEN_979; // @[AxiStoreQueue.scala 166:35:@1787.4]
  wire  _T_3603; // @[AxiStoreQueue.scala 168:54:@1800.6]
  wire  _T_3604; // @[AxiStoreQueue.scala 168:36:@1801.6]
  wire  _GEN_980; // @[AxiStoreQueue.scala 168:75:@1802.6]
  wire  _GEN_981; // @[AxiStoreQueue.scala 166:35:@1796.4]
  wire  _T_3608; // @[AxiStoreQueue.scala 168:54:@1809.6]
  wire  _T_3609; // @[AxiStoreQueue.scala 168:36:@1810.6]
  wire  _GEN_982; // @[AxiStoreQueue.scala 168:75:@1811.6]
  wire  _GEN_983; // @[AxiStoreQueue.scala 166:35:@1805.4]
  wire  _T_3613; // @[AxiStoreQueue.scala 168:54:@1818.6]
  wire  _T_3614; // @[AxiStoreQueue.scala 168:36:@1819.6]
  wire  _GEN_984; // @[AxiStoreQueue.scala 168:75:@1820.6]
  wire  _GEN_985; // @[AxiStoreQueue.scala 166:35:@1814.4]
  wire  _T_3618; // @[AxiStoreQueue.scala 168:54:@1827.6]
  wire  _T_3619; // @[AxiStoreQueue.scala 168:36:@1828.6]
  wire  _GEN_986; // @[AxiStoreQueue.scala 168:75:@1829.6]
  wire  _GEN_987; // @[AxiStoreQueue.scala 166:35:@1823.4]
  wire  _T_3623; // @[AxiStoreQueue.scala 168:54:@1836.6]
  wire  _T_3624; // @[AxiStoreQueue.scala 168:36:@1837.6]
  wire  _GEN_988; // @[AxiStoreQueue.scala 168:75:@1838.6]
  wire  _GEN_989; // @[AxiStoreQueue.scala 166:35:@1832.4]
  wire  _T_3628; // @[AxiStoreQueue.scala 168:54:@1845.6]
  wire  _T_3629; // @[AxiStoreQueue.scala 168:36:@1846.6]
  wire  _GEN_990; // @[AxiStoreQueue.scala 168:75:@1847.6]
  wire  _GEN_991; // @[AxiStoreQueue.scala 166:35:@1841.4]
  wire  entriesPorts_0_0; // @[AxiStoreQueue.scala 185:72:@1851.4]
  wire  entriesPorts_0_1; // @[AxiStoreQueue.scala 185:72:@1853.4]
  wire  entriesPorts_0_2; // @[AxiStoreQueue.scala 185:72:@1855.4]
  wire  entriesPorts_0_3; // @[AxiStoreQueue.scala 185:72:@1857.4]
  wire  entriesPorts_0_4; // @[AxiStoreQueue.scala 185:72:@1859.4]
  wire  entriesPorts_0_5; // @[AxiStoreQueue.scala 185:72:@1861.4]
  wire  entriesPorts_0_6; // @[AxiStoreQueue.scala 185:72:@1863.4]
  wire  entriesPorts_0_7; // @[AxiStoreQueue.scala 185:72:@1865.4]
  wire  entriesPorts_0_8; // @[AxiStoreQueue.scala 185:72:@1867.4]
  wire  entriesPorts_0_9; // @[AxiStoreQueue.scala 185:72:@1869.4]
  wire  entriesPorts_0_10; // @[AxiStoreQueue.scala 185:72:@1871.4]
  wire  entriesPorts_0_11; // @[AxiStoreQueue.scala 185:72:@1873.4]
  wire  entriesPorts_0_12; // @[AxiStoreQueue.scala 185:72:@1875.4]
  wire  entriesPorts_0_13; // @[AxiStoreQueue.scala 185:72:@1877.4]
  wire  entriesPorts_0_14; // @[AxiStoreQueue.scala 185:72:@1879.4]
  wire  entriesPorts_0_15; // @[AxiStoreQueue.scala 185:72:@1881.4]
  wire  _T_4114; // @[AxiStoreQueue.scala 197:91:@1885.4]
  wire  _T_4115; // @[AxiStoreQueue.scala 197:88:@1886.4]
  wire  _T_4117; // @[AxiStoreQueue.scala 197:91:@1887.4]
  wire  _T_4118; // @[AxiStoreQueue.scala 197:88:@1888.4]
  wire  _T_4120; // @[AxiStoreQueue.scala 197:91:@1889.4]
  wire  _T_4121; // @[AxiStoreQueue.scala 197:88:@1890.4]
  wire  _T_4123; // @[AxiStoreQueue.scala 197:91:@1891.4]
  wire  _T_4124; // @[AxiStoreQueue.scala 197:88:@1892.4]
  wire  _T_4126; // @[AxiStoreQueue.scala 197:91:@1893.4]
  wire  _T_4127; // @[AxiStoreQueue.scala 197:88:@1894.4]
  wire  _T_4129; // @[AxiStoreQueue.scala 197:91:@1895.4]
  wire  _T_4130; // @[AxiStoreQueue.scala 197:88:@1896.4]
  wire  _T_4132; // @[AxiStoreQueue.scala 197:91:@1897.4]
  wire  _T_4133; // @[AxiStoreQueue.scala 197:88:@1898.4]
  wire  _T_4135; // @[AxiStoreQueue.scala 197:91:@1899.4]
  wire  _T_4136; // @[AxiStoreQueue.scala 197:88:@1900.4]
  wire  _T_4138; // @[AxiStoreQueue.scala 197:91:@1901.4]
  wire  _T_4139; // @[AxiStoreQueue.scala 197:88:@1902.4]
  wire  _T_4141; // @[AxiStoreQueue.scala 197:91:@1903.4]
  wire  _T_4142; // @[AxiStoreQueue.scala 197:88:@1904.4]
  wire  _T_4144; // @[AxiStoreQueue.scala 197:91:@1905.4]
  wire  _T_4145; // @[AxiStoreQueue.scala 197:88:@1906.4]
  wire  _T_4147; // @[AxiStoreQueue.scala 197:91:@1907.4]
  wire  _T_4148; // @[AxiStoreQueue.scala 197:88:@1908.4]
  wire  _T_4150; // @[AxiStoreQueue.scala 197:91:@1909.4]
  wire  _T_4151; // @[AxiStoreQueue.scala 197:88:@1910.4]
  wire  _T_4153; // @[AxiStoreQueue.scala 197:91:@1911.4]
  wire  _T_4154; // @[AxiStoreQueue.scala 197:88:@1912.4]
  wire  _T_4156; // @[AxiStoreQueue.scala 197:91:@1913.4]
  wire  _T_4157; // @[AxiStoreQueue.scala 197:88:@1914.4]
  wire  _T_4159; // @[AxiStoreQueue.scala 197:91:@1915.4]
  wire  _T_4160; // @[AxiStoreQueue.scala 197:88:@1916.4]
  wire  _T_4184; // @[AxiStoreQueue.scala 198:91:@1934.4]
  wire  _T_4185; // @[AxiStoreQueue.scala 198:88:@1935.4]
  wire  _T_4187; // @[AxiStoreQueue.scala 198:91:@1936.4]
  wire  _T_4188; // @[AxiStoreQueue.scala 198:88:@1937.4]
  wire  _T_4190; // @[AxiStoreQueue.scala 198:91:@1938.4]
  wire  _T_4191; // @[AxiStoreQueue.scala 198:88:@1939.4]
  wire  _T_4193; // @[AxiStoreQueue.scala 198:91:@1940.4]
  wire  _T_4194; // @[AxiStoreQueue.scala 198:88:@1941.4]
  wire  _T_4196; // @[AxiStoreQueue.scala 198:91:@1942.4]
  wire  _T_4197; // @[AxiStoreQueue.scala 198:88:@1943.4]
  wire  _T_4199; // @[AxiStoreQueue.scala 198:91:@1944.4]
  wire  _T_4200; // @[AxiStoreQueue.scala 198:88:@1945.4]
  wire  _T_4202; // @[AxiStoreQueue.scala 198:91:@1946.4]
  wire  _T_4203; // @[AxiStoreQueue.scala 198:88:@1947.4]
  wire  _T_4205; // @[AxiStoreQueue.scala 198:91:@1948.4]
  wire  _T_4206; // @[AxiStoreQueue.scala 198:88:@1949.4]
  wire  _T_4208; // @[AxiStoreQueue.scala 198:91:@1950.4]
  wire  _T_4209; // @[AxiStoreQueue.scala 198:88:@1951.4]
  wire  _T_4211; // @[AxiStoreQueue.scala 198:91:@1952.4]
  wire  _T_4212; // @[AxiStoreQueue.scala 198:88:@1953.4]
  wire  _T_4214; // @[AxiStoreQueue.scala 198:91:@1954.4]
  wire  _T_4215; // @[AxiStoreQueue.scala 198:88:@1955.4]
  wire  _T_4217; // @[AxiStoreQueue.scala 198:91:@1956.4]
  wire  _T_4218; // @[AxiStoreQueue.scala 198:88:@1957.4]
  wire  _T_4220; // @[AxiStoreQueue.scala 198:91:@1958.4]
  wire  _T_4221; // @[AxiStoreQueue.scala 198:88:@1959.4]
  wire  _T_4223; // @[AxiStoreQueue.scala 198:91:@1960.4]
  wire  _T_4224; // @[AxiStoreQueue.scala 198:88:@1961.4]
  wire  _T_4226; // @[AxiStoreQueue.scala 198:91:@1962.4]
  wire  _T_4227; // @[AxiStoreQueue.scala 198:88:@1963.4]
  wire  _T_4229; // @[AxiStoreQueue.scala 198:91:@1964.4]
  wire  _T_4230; // @[AxiStoreQueue.scala 198:88:@1965.4]
  wire [15:0] _T_4255; // @[OneHot.scala 52:12:@1984.4]
  wire  _T_4257; // @[util.scala 33:60:@1986.4]
  wire  _T_4258; // @[util.scala 33:60:@1987.4]
  wire  _T_4259; // @[util.scala 33:60:@1988.4]
  wire  _T_4260; // @[util.scala 33:60:@1989.4]
  wire  _T_4261; // @[util.scala 33:60:@1990.4]
  wire  _T_4262; // @[util.scala 33:60:@1991.4]
  wire  _T_4263; // @[util.scala 33:60:@1992.4]
  wire  _T_4264; // @[util.scala 33:60:@1993.4]
  wire  _T_4265; // @[util.scala 33:60:@1994.4]
  wire  _T_4266; // @[util.scala 33:60:@1995.4]
  wire  _T_4267; // @[util.scala 33:60:@1996.4]
  wire  _T_4268; // @[util.scala 33:60:@1997.4]
  wire  _T_4269; // @[util.scala 33:60:@1998.4]
  wire  _T_4270; // @[util.scala 33:60:@1999.4]
  wire  _T_4271; // @[util.scala 33:60:@2000.4]
  wire  _T_4272; // @[util.scala 33:60:@2001.4]
  wire [15:0] _T_4313; // @[Mux.scala 31:69:@2019.4]
  wire [15:0] _T_4314; // @[Mux.scala 31:69:@2020.4]
  wire [15:0] _T_4315; // @[Mux.scala 31:69:@2021.4]
  wire [15:0] _T_4316; // @[Mux.scala 31:69:@2022.4]
  wire [15:0] _T_4317; // @[Mux.scala 31:69:@2023.4]
  wire [15:0] _T_4318; // @[Mux.scala 31:69:@2024.4]
  wire [15:0] _T_4319; // @[Mux.scala 31:69:@2025.4]
  wire [15:0] _T_4320; // @[Mux.scala 31:69:@2026.4]
  wire [15:0] _T_4321; // @[Mux.scala 31:69:@2027.4]
  wire [15:0] _T_4322; // @[Mux.scala 31:69:@2028.4]
  wire [15:0] _T_4323; // @[Mux.scala 31:69:@2029.4]
  wire [15:0] _T_4324; // @[Mux.scala 31:69:@2030.4]
  wire [15:0] _T_4325; // @[Mux.scala 31:69:@2031.4]
  wire [15:0] _T_4326; // @[Mux.scala 31:69:@2032.4]
  wire [15:0] _T_4327; // @[Mux.scala 31:69:@2033.4]
  wire [15:0] _T_4328; // @[Mux.scala 31:69:@2034.4]
  wire  _T_4329; // @[OneHot.scala 66:30:@2035.4]
  wire  _T_4330; // @[OneHot.scala 66:30:@2036.4]
  wire  _T_4331; // @[OneHot.scala 66:30:@2037.4]
  wire  _T_4332; // @[OneHot.scala 66:30:@2038.4]
  wire  _T_4333; // @[OneHot.scala 66:30:@2039.4]
  wire  _T_4334; // @[OneHot.scala 66:30:@2040.4]
  wire  _T_4335; // @[OneHot.scala 66:30:@2041.4]
  wire  _T_4336; // @[OneHot.scala 66:30:@2042.4]
  wire  _T_4337; // @[OneHot.scala 66:30:@2043.4]
  wire  _T_4338; // @[OneHot.scala 66:30:@2044.4]
  wire  _T_4339; // @[OneHot.scala 66:30:@2045.4]
  wire  _T_4340; // @[OneHot.scala 66:30:@2046.4]
  wire  _T_4341; // @[OneHot.scala 66:30:@2047.4]
  wire  _T_4342; // @[OneHot.scala 66:30:@2048.4]
  wire  _T_4343; // @[OneHot.scala 66:30:@2049.4]
  wire  _T_4344; // @[OneHot.scala 66:30:@2050.4]
  wire [15:0] _T_4385; // @[Mux.scala 31:69:@2068.4]
  wire [15:0] _T_4386; // @[Mux.scala 31:69:@2069.4]
  wire [15:0] _T_4387; // @[Mux.scala 31:69:@2070.4]
  wire [15:0] _T_4388; // @[Mux.scala 31:69:@2071.4]
  wire [15:0] _T_4389; // @[Mux.scala 31:69:@2072.4]
  wire [15:0] _T_4390; // @[Mux.scala 31:69:@2073.4]
  wire [15:0] _T_4391; // @[Mux.scala 31:69:@2074.4]
  wire [15:0] _T_4392; // @[Mux.scala 31:69:@2075.4]
  wire [15:0] _T_4393; // @[Mux.scala 31:69:@2076.4]
  wire [15:0] _T_4394; // @[Mux.scala 31:69:@2077.4]
  wire [15:0] _T_4395; // @[Mux.scala 31:69:@2078.4]
  wire [15:0] _T_4396; // @[Mux.scala 31:69:@2079.4]
  wire [15:0] _T_4397; // @[Mux.scala 31:69:@2080.4]
  wire [15:0] _T_4398; // @[Mux.scala 31:69:@2081.4]
  wire [15:0] _T_4399; // @[Mux.scala 31:69:@2082.4]
  wire [15:0] _T_4400; // @[Mux.scala 31:69:@2083.4]
  wire  _T_4401; // @[OneHot.scala 66:30:@2084.4]
  wire  _T_4402; // @[OneHot.scala 66:30:@2085.4]
  wire  _T_4403; // @[OneHot.scala 66:30:@2086.4]
  wire  _T_4404; // @[OneHot.scala 66:30:@2087.4]
  wire  _T_4405; // @[OneHot.scala 66:30:@2088.4]
  wire  _T_4406; // @[OneHot.scala 66:30:@2089.4]
  wire  _T_4407; // @[OneHot.scala 66:30:@2090.4]
  wire  _T_4408; // @[OneHot.scala 66:30:@2091.4]
  wire  _T_4409; // @[OneHot.scala 66:30:@2092.4]
  wire  _T_4410; // @[OneHot.scala 66:30:@2093.4]
  wire  _T_4411; // @[OneHot.scala 66:30:@2094.4]
  wire  _T_4412; // @[OneHot.scala 66:30:@2095.4]
  wire  _T_4413; // @[OneHot.scala 66:30:@2096.4]
  wire  _T_4414; // @[OneHot.scala 66:30:@2097.4]
  wire  _T_4415; // @[OneHot.scala 66:30:@2098.4]
  wire  _T_4416; // @[OneHot.scala 66:30:@2099.4]
  wire [15:0] _T_4457; // @[Mux.scala 31:69:@2117.4]
  wire [15:0] _T_4458; // @[Mux.scala 31:69:@2118.4]
  wire [15:0] _T_4459; // @[Mux.scala 31:69:@2119.4]
  wire [15:0] _T_4460; // @[Mux.scala 31:69:@2120.4]
  wire [15:0] _T_4461; // @[Mux.scala 31:69:@2121.4]
  wire [15:0] _T_4462; // @[Mux.scala 31:69:@2122.4]
  wire [15:0] _T_4463; // @[Mux.scala 31:69:@2123.4]
  wire [15:0] _T_4464; // @[Mux.scala 31:69:@2124.4]
  wire [15:0] _T_4465; // @[Mux.scala 31:69:@2125.4]
  wire [15:0] _T_4466; // @[Mux.scala 31:69:@2126.4]
  wire [15:0] _T_4467; // @[Mux.scala 31:69:@2127.4]
  wire [15:0] _T_4468; // @[Mux.scala 31:69:@2128.4]
  wire [15:0] _T_4469; // @[Mux.scala 31:69:@2129.4]
  wire [15:0] _T_4470; // @[Mux.scala 31:69:@2130.4]
  wire [15:0] _T_4471; // @[Mux.scala 31:69:@2131.4]
  wire [15:0] _T_4472; // @[Mux.scala 31:69:@2132.4]
  wire  _T_4473; // @[OneHot.scala 66:30:@2133.4]
  wire  _T_4474; // @[OneHot.scala 66:30:@2134.4]
  wire  _T_4475; // @[OneHot.scala 66:30:@2135.4]
  wire  _T_4476; // @[OneHot.scala 66:30:@2136.4]
  wire  _T_4477; // @[OneHot.scala 66:30:@2137.4]
  wire  _T_4478; // @[OneHot.scala 66:30:@2138.4]
  wire  _T_4479; // @[OneHot.scala 66:30:@2139.4]
  wire  _T_4480; // @[OneHot.scala 66:30:@2140.4]
  wire  _T_4481; // @[OneHot.scala 66:30:@2141.4]
  wire  _T_4482; // @[OneHot.scala 66:30:@2142.4]
  wire  _T_4483; // @[OneHot.scala 66:30:@2143.4]
  wire  _T_4484; // @[OneHot.scala 66:30:@2144.4]
  wire  _T_4485; // @[OneHot.scala 66:30:@2145.4]
  wire  _T_4486; // @[OneHot.scala 66:30:@2146.4]
  wire  _T_4487; // @[OneHot.scala 66:30:@2147.4]
  wire  _T_4488; // @[OneHot.scala 66:30:@2148.4]
  wire [15:0] _T_4529; // @[Mux.scala 31:69:@2166.4]
  wire [15:0] _T_4530; // @[Mux.scala 31:69:@2167.4]
  wire [15:0] _T_4531; // @[Mux.scala 31:69:@2168.4]
  wire [15:0] _T_4532; // @[Mux.scala 31:69:@2169.4]
  wire [15:0] _T_4533; // @[Mux.scala 31:69:@2170.4]
  wire [15:0] _T_4534; // @[Mux.scala 31:69:@2171.4]
  wire [15:0] _T_4535; // @[Mux.scala 31:69:@2172.4]
  wire [15:0] _T_4536; // @[Mux.scala 31:69:@2173.4]
  wire [15:0] _T_4537; // @[Mux.scala 31:69:@2174.4]
  wire [15:0] _T_4538; // @[Mux.scala 31:69:@2175.4]
  wire [15:0] _T_4539; // @[Mux.scala 31:69:@2176.4]
  wire [15:0] _T_4540; // @[Mux.scala 31:69:@2177.4]
  wire [15:0] _T_4541; // @[Mux.scala 31:69:@2178.4]
  wire [15:0] _T_4542; // @[Mux.scala 31:69:@2179.4]
  wire [15:0] _T_4543; // @[Mux.scala 31:69:@2180.4]
  wire [15:0] _T_4544; // @[Mux.scala 31:69:@2181.4]
  wire  _T_4545; // @[OneHot.scala 66:30:@2182.4]
  wire  _T_4546; // @[OneHot.scala 66:30:@2183.4]
  wire  _T_4547; // @[OneHot.scala 66:30:@2184.4]
  wire  _T_4548; // @[OneHot.scala 66:30:@2185.4]
  wire  _T_4549; // @[OneHot.scala 66:30:@2186.4]
  wire  _T_4550; // @[OneHot.scala 66:30:@2187.4]
  wire  _T_4551; // @[OneHot.scala 66:30:@2188.4]
  wire  _T_4552; // @[OneHot.scala 66:30:@2189.4]
  wire  _T_4553; // @[OneHot.scala 66:30:@2190.4]
  wire  _T_4554; // @[OneHot.scala 66:30:@2191.4]
  wire  _T_4555; // @[OneHot.scala 66:30:@2192.4]
  wire  _T_4556; // @[OneHot.scala 66:30:@2193.4]
  wire  _T_4557; // @[OneHot.scala 66:30:@2194.4]
  wire  _T_4558; // @[OneHot.scala 66:30:@2195.4]
  wire  _T_4559; // @[OneHot.scala 66:30:@2196.4]
  wire  _T_4560; // @[OneHot.scala 66:30:@2197.4]
  wire [15:0] _T_4601; // @[Mux.scala 31:69:@2215.4]
  wire [15:0] _T_4602; // @[Mux.scala 31:69:@2216.4]
  wire [15:0] _T_4603; // @[Mux.scala 31:69:@2217.4]
  wire [15:0] _T_4604; // @[Mux.scala 31:69:@2218.4]
  wire [15:0] _T_4605; // @[Mux.scala 31:69:@2219.4]
  wire [15:0] _T_4606; // @[Mux.scala 31:69:@2220.4]
  wire [15:0] _T_4607; // @[Mux.scala 31:69:@2221.4]
  wire [15:0] _T_4608; // @[Mux.scala 31:69:@2222.4]
  wire [15:0] _T_4609; // @[Mux.scala 31:69:@2223.4]
  wire [15:0] _T_4610; // @[Mux.scala 31:69:@2224.4]
  wire [15:0] _T_4611; // @[Mux.scala 31:69:@2225.4]
  wire [15:0] _T_4612; // @[Mux.scala 31:69:@2226.4]
  wire [15:0] _T_4613; // @[Mux.scala 31:69:@2227.4]
  wire [15:0] _T_4614; // @[Mux.scala 31:69:@2228.4]
  wire [15:0] _T_4615; // @[Mux.scala 31:69:@2229.4]
  wire [15:0] _T_4616; // @[Mux.scala 31:69:@2230.4]
  wire  _T_4617; // @[OneHot.scala 66:30:@2231.4]
  wire  _T_4618; // @[OneHot.scala 66:30:@2232.4]
  wire  _T_4619; // @[OneHot.scala 66:30:@2233.4]
  wire  _T_4620; // @[OneHot.scala 66:30:@2234.4]
  wire  _T_4621; // @[OneHot.scala 66:30:@2235.4]
  wire  _T_4622; // @[OneHot.scala 66:30:@2236.4]
  wire  _T_4623; // @[OneHot.scala 66:30:@2237.4]
  wire  _T_4624; // @[OneHot.scala 66:30:@2238.4]
  wire  _T_4625; // @[OneHot.scala 66:30:@2239.4]
  wire  _T_4626; // @[OneHot.scala 66:30:@2240.4]
  wire  _T_4627; // @[OneHot.scala 66:30:@2241.4]
  wire  _T_4628; // @[OneHot.scala 66:30:@2242.4]
  wire  _T_4629; // @[OneHot.scala 66:30:@2243.4]
  wire  _T_4630; // @[OneHot.scala 66:30:@2244.4]
  wire  _T_4631; // @[OneHot.scala 66:30:@2245.4]
  wire  _T_4632; // @[OneHot.scala 66:30:@2246.4]
  wire [15:0] _T_4673; // @[Mux.scala 31:69:@2264.4]
  wire [15:0] _T_4674; // @[Mux.scala 31:69:@2265.4]
  wire [15:0] _T_4675; // @[Mux.scala 31:69:@2266.4]
  wire [15:0] _T_4676; // @[Mux.scala 31:69:@2267.4]
  wire [15:0] _T_4677; // @[Mux.scala 31:69:@2268.4]
  wire [15:0] _T_4678; // @[Mux.scala 31:69:@2269.4]
  wire [15:0] _T_4679; // @[Mux.scala 31:69:@2270.4]
  wire [15:0] _T_4680; // @[Mux.scala 31:69:@2271.4]
  wire [15:0] _T_4681; // @[Mux.scala 31:69:@2272.4]
  wire [15:0] _T_4682; // @[Mux.scala 31:69:@2273.4]
  wire [15:0] _T_4683; // @[Mux.scala 31:69:@2274.4]
  wire [15:0] _T_4684; // @[Mux.scala 31:69:@2275.4]
  wire [15:0] _T_4685; // @[Mux.scala 31:69:@2276.4]
  wire [15:0] _T_4686; // @[Mux.scala 31:69:@2277.4]
  wire [15:0] _T_4687; // @[Mux.scala 31:69:@2278.4]
  wire [15:0] _T_4688; // @[Mux.scala 31:69:@2279.4]
  wire  _T_4689; // @[OneHot.scala 66:30:@2280.4]
  wire  _T_4690; // @[OneHot.scala 66:30:@2281.4]
  wire  _T_4691; // @[OneHot.scala 66:30:@2282.4]
  wire  _T_4692; // @[OneHot.scala 66:30:@2283.4]
  wire  _T_4693; // @[OneHot.scala 66:30:@2284.4]
  wire  _T_4694; // @[OneHot.scala 66:30:@2285.4]
  wire  _T_4695; // @[OneHot.scala 66:30:@2286.4]
  wire  _T_4696; // @[OneHot.scala 66:30:@2287.4]
  wire  _T_4697; // @[OneHot.scala 66:30:@2288.4]
  wire  _T_4698; // @[OneHot.scala 66:30:@2289.4]
  wire  _T_4699; // @[OneHot.scala 66:30:@2290.4]
  wire  _T_4700; // @[OneHot.scala 66:30:@2291.4]
  wire  _T_4701; // @[OneHot.scala 66:30:@2292.4]
  wire  _T_4702; // @[OneHot.scala 66:30:@2293.4]
  wire  _T_4703; // @[OneHot.scala 66:30:@2294.4]
  wire  _T_4704; // @[OneHot.scala 66:30:@2295.4]
  wire [15:0] _T_4745; // @[Mux.scala 31:69:@2313.4]
  wire [15:0] _T_4746; // @[Mux.scala 31:69:@2314.4]
  wire [15:0] _T_4747; // @[Mux.scala 31:69:@2315.4]
  wire [15:0] _T_4748; // @[Mux.scala 31:69:@2316.4]
  wire [15:0] _T_4749; // @[Mux.scala 31:69:@2317.4]
  wire [15:0] _T_4750; // @[Mux.scala 31:69:@2318.4]
  wire [15:0] _T_4751; // @[Mux.scala 31:69:@2319.4]
  wire [15:0] _T_4752; // @[Mux.scala 31:69:@2320.4]
  wire [15:0] _T_4753; // @[Mux.scala 31:69:@2321.4]
  wire [15:0] _T_4754; // @[Mux.scala 31:69:@2322.4]
  wire [15:0] _T_4755; // @[Mux.scala 31:69:@2323.4]
  wire [15:0] _T_4756; // @[Mux.scala 31:69:@2324.4]
  wire [15:0] _T_4757; // @[Mux.scala 31:69:@2325.4]
  wire [15:0] _T_4758; // @[Mux.scala 31:69:@2326.4]
  wire [15:0] _T_4759; // @[Mux.scala 31:69:@2327.4]
  wire [15:0] _T_4760; // @[Mux.scala 31:69:@2328.4]
  wire  _T_4761; // @[OneHot.scala 66:30:@2329.4]
  wire  _T_4762; // @[OneHot.scala 66:30:@2330.4]
  wire  _T_4763; // @[OneHot.scala 66:30:@2331.4]
  wire  _T_4764; // @[OneHot.scala 66:30:@2332.4]
  wire  _T_4765; // @[OneHot.scala 66:30:@2333.4]
  wire  _T_4766; // @[OneHot.scala 66:30:@2334.4]
  wire  _T_4767; // @[OneHot.scala 66:30:@2335.4]
  wire  _T_4768; // @[OneHot.scala 66:30:@2336.4]
  wire  _T_4769; // @[OneHot.scala 66:30:@2337.4]
  wire  _T_4770; // @[OneHot.scala 66:30:@2338.4]
  wire  _T_4771; // @[OneHot.scala 66:30:@2339.4]
  wire  _T_4772; // @[OneHot.scala 66:30:@2340.4]
  wire  _T_4773; // @[OneHot.scala 66:30:@2341.4]
  wire  _T_4774; // @[OneHot.scala 66:30:@2342.4]
  wire  _T_4775; // @[OneHot.scala 66:30:@2343.4]
  wire  _T_4776; // @[OneHot.scala 66:30:@2344.4]
  wire [15:0] _T_4817; // @[Mux.scala 31:69:@2362.4]
  wire [15:0] _T_4818; // @[Mux.scala 31:69:@2363.4]
  wire [15:0] _T_4819; // @[Mux.scala 31:69:@2364.4]
  wire [15:0] _T_4820; // @[Mux.scala 31:69:@2365.4]
  wire [15:0] _T_4821; // @[Mux.scala 31:69:@2366.4]
  wire [15:0] _T_4822; // @[Mux.scala 31:69:@2367.4]
  wire [15:0] _T_4823; // @[Mux.scala 31:69:@2368.4]
  wire [15:0] _T_4824; // @[Mux.scala 31:69:@2369.4]
  wire [15:0] _T_4825; // @[Mux.scala 31:69:@2370.4]
  wire [15:0] _T_4826; // @[Mux.scala 31:69:@2371.4]
  wire [15:0] _T_4827; // @[Mux.scala 31:69:@2372.4]
  wire [15:0] _T_4828; // @[Mux.scala 31:69:@2373.4]
  wire [15:0] _T_4829; // @[Mux.scala 31:69:@2374.4]
  wire [15:0] _T_4830; // @[Mux.scala 31:69:@2375.4]
  wire [15:0] _T_4831; // @[Mux.scala 31:69:@2376.4]
  wire [15:0] _T_4832; // @[Mux.scala 31:69:@2377.4]
  wire  _T_4833; // @[OneHot.scala 66:30:@2378.4]
  wire  _T_4834; // @[OneHot.scala 66:30:@2379.4]
  wire  _T_4835; // @[OneHot.scala 66:30:@2380.4]
  wire  _T_4836; // @[OneHot.scala 66:30:@2381.4]
  wire  _T_4837; // @[OneHot.scala 66:30:@2382.4]
  wire  _T_4838; // @[OneHot.scala 66:30:@2383.4]
  wire  _T_4839; // @[OneHot.scala 66:30:@2384.4]
  wire  _T_4840; // @[OneHot.scala 66:30:@2385.4]
  wire  _T_4841; // @[OneHot.scala 66:30:@2386.4]
  wire  _T_4842; // @[OneHot.scala 66:30:@2387.4]
  wire  _T_4843; // @[OneHot.scala 66:30:@2388.4]
  wire  _T_4844; // @[OneHot.scala 66:30:@2389.4]
  wire  _T_4845; // @[OneHot.scala 66:30:@2390.4]
  wire  _T_4846; // @[OneHot.scala 66:30:@2391.4]
  wire  _T_4847; // @[OneHot.scala 66:30:@2392.4]
  wire  _T_4848; // @[OneHot.scala 66:30:@2393.4]
  wire [15:0] _T_4889; // @[Mux.scala 31:69:@2411.4]
  wire [15:0] _T_4890; // @[Mux.scala 31:69:@2412.4]
  wire [15:0] _T_4891; // @[Mux.scala 31:69:@2413.4]
  wire [15:0] _T_4892; // @[Mux.scala 31:69:@2414.4]
  wire [15:0] _T_4893; // @[Mux.scala 31:69:@2415.4]
  wire [15:0] _T_4894; // @[Mux.scala 31:69:@2416.4]
  wire [15:0] _T_4895; // @[Mux.scala 31:69:@2417.4]
  wire [15:0] _T_4896; // @[Mux.scala 31:69:@2418.4]
  wire [15:0] _T_4897; // @[Mux.scala 31:69:@2419.4]
  wire [15:0] _T_4898; // @[Mux.scala 31:69:@2420.4]
  wire [15:0] _T_4899; // @[Mux.scala 31:69:@2421.4]
  wire [15:0] _T_4900; // @[Mux.scala 31:69:@2422.4]
  wire [15:0] _T_4901; // @[Mux.scala 31:69:@2423.4]
  wire [15:0] _T_4902; // @[Mux.scala 31:69:@2424.4]
  wire [15:0] _T_4903; // @[Mux.scala 31:69:@2425.4]
  wire [15:0] _T_4904; // @[Mux.scala 31:69:@2426.4]
  wire  _T_4905; // @[OneHot.scala 66:30:@2427.4]
  wire  _T_4906; // @[OneHot.scala 66:30:@2428.4]
  wire  _T_4907; // @[OneHot.scala 66:30:@2429.4]
  wire  _T_4908; // @[OneHot.scala 66:30:@2430.4]
  wire  _T_4909; // @[OneHot.scala 66:30:@2431.4]
  wire  _T_4910; // @[OneHot.scala 66:30:@2432.4]
  wire  _T_4911; // @[OneHot.scala 66:30:@2433.4]
  wire  _T_4912; // @[OneHot.scala 66:30:@2434.4]
  wire  _T_4913; // @[OneHot.scala 66:30:@2435.4]
  wire  _T_4914; // @[OneHot.scala 66:30:@2436.4]
  wire  _T_4915; // @[OneHot.scala 66:30:@2437.4]
  wire  _T_4916; // @[OneHot.scala 66:30:@2438.4]
  wire  _T_4917; // @[OneHot.scala 66:30:@2439.4]
  wire  _T_4918; // @[OneHot.scala 66:30:@2440.4]
  wire  _T_4919; // @[OneHot.scala 66:30:@2441.4]
  wire  _T_4920; // @[OneHot.scala 66:30:@2442.4]
  wire [15:0] _T_4961; // @[Mux.scala 31:69:@2460.4]
  wire [15:0] _T_4962; // @[Mux.scala 31:69:@2461.4]
  wire [15:0] _T_4963; // @[Mux.scala 31:69:@2462.4]
  wire [15:0] _T_4964; // @[Mux.scala 31:69:@2463.4]
  wire [15:0] _T_4965; // @[Mux.scala 31:69:@2464.4]
  wire [15:0] _T_4966; // @[Mux.scala 31:69:@2465.4]
  wire [15:0] _T_4967; // @[Mux.scala 31:69:@2466.4]
  wire [15:0] _T_4968; // @[Mux.scala 31:69:@2467.4]
  wire [15:0] _T_4969; // @[Mux.scala 31:69:@2468.4]
  wire [15:0] _T_4970; // @[Mux.scala 31:69:@2469.4]
  wire [15:0] _T_4971; // @[Mux.scala 31:69:@2470.4]
  wire [15:0] _T_4972; // @[Mux.scala 31:69:@2471.4]
  wire [15:0] _T_4973; // @[Mux.scala 31:69:@2472.4]
  wire [15:0] _T_4974; // @[Mux.scala 31:69:@2473.4]
  wire [15:0] _T_4975; // @[Mux.scala 31:69:@2474.4]
  wire [15:0] _T_4976; // @[Mux.scala 31:69:@2475.4]
  wire  _T_4977; // @[OneHot.scala 66:30:@2476.4]
  wire  _T_4978; // @[OneHot.scala 66:30:@2477.4]
  wire  _T_4979; // @[OneHot.scala 66:30:@2478.4]
  wire  _T_4980; // @[OneHot.scala 66:30:@2479.4]
  wire  _T_4981; // @[OneHot.scala 66:30:@2480.4]
  wire  _T_4982; // @[OneHot.scala 66:30:@2481.4]
  wire  _T_4983; // @[OneHot.scala 66:30:@2482.4]
  wire  _T_4984; // @[OneHot.scala 66:30:@2483.4]
  wire  _T_4985; // @[OneHot.scala 66:30:@2484.4]
  wire  _T_4986; // @[OneHot.scala 66:30:@2485.4]
  wire  _T_4987; // @[OneHot.scala 66:30:@2486.4]
  wire  _T_4988; // @[OneHot.scala 66:30:@2487.4]
  wire  _T_4989; // @[OneHot.scala 66:30:@2488.4]
  wire  _T_4990; // @[OneHot.scala 66:30:@2489.4]
  wire  _T_4991; // @[OneHot.scala 66:30:@2490.4]
  wire  _T_4992; // @[OneHot.scala 66:30:@2491.4]
  wire [15:0] _T_5033; // @[Mux.scala 31:69:@2509.4]
  wire [15:0] _T_5034; // @[Mux.scala 31:69:@2510.4]
  wire [15:0] _T_5035; // @[Mux.scala 31:69:@2511.4]
  wire [15:0] _T_5036; // @[Mux.scala 31:69:@2512.4]
  wire [15:0] _T_5037; // @[Mux.scala 31:69:@2513.4]
  wire [15:0] _T_5038; // @[Mux.scala 31:69:@2514.4]
  wire [15:0] _T_5039; // @[Mux.scala 31:69:@2515.4]
  wire [15:0] _T_5040; // @[Mux.scala 31:69:@2516.4]
  wire [15:0] _T_5041; // @[Mux.scala 31:69:@2517.4]
  wire [15:0] _T_5042; // @[Mux.scala 31:69:@2518.4]
  wire [15:0] _T_5043; // @[Mux.scala 31:69:@2519.4]
  wire [15:0] _T_5044; // @[Mux.scala 31:69:@2520.4]
  wire [15:0] _T_5045; // @[Mux.scala 31:69:@2521.4]
  wire [15:0] _T_5046; // @[Mux.scala 31:69:@2522.4]
  wire [15:0] _T_5047; // @[Mux.scala 31:69:@2523.4]
  wire [15:0] _T_5048; // @[Mux.scala 31:69:@2524.4]
  wire  _T_5049; // @[OneHot.scala 66:30:@2525.4]
  wire  _T_5050; // @[OneHot.scala 66:30:@2526.4]
  wire  _T_5051; // @[OneHot.scala 66:30:@2527.4]
  wire  _T_5052; // @[OneHot.scala 66:30:@2528.4]
  wire  _T_5053; // @[OneHot.scala 66:30:@2529.4]
  wire  _T_5054; // @[OneHot.scala 66:30:@2530.4]
  wire  _T_5055; // @[OneHot.scala 66:30:@2531.4]
  wire  _T_5056; // @[OneHot.scala 66:30:@2532.4]
  wire  _T_5057; // @[OneHot.scala 66:30:@2533.4]
  wire  _T_5058; // @[OneHot.scala 66:30:@2534.4]
  wire  _T_5059; // @[OneHot.scala 66:30:@2535.4]
  wire  _T_5060; // @[OneHot.scala 66:30:@2536.4]
  wire  _T_5061; // @[OneHot.scala 66:30:@2537.4]
  wire  _T_5062; // @[OneHot.scala 66:30:@2538.4]
  wire  _T_5063; // @[OneHot.scala 66:30:@2539.4]
  wire  _T_5064; // @[OneHot.scala 66:30:@2540.4]
  wire [15:0] _T_5105; // @[Mux.scala 31:69:@2558.4]
  wire [15:0] _T_5106; // @[Mux.scala 31:69:@2559.4]
  wire [15:0] _T_5107; // @[Mux.scala 31:69:@2560.4]
  wire [15:0] _T_5108; // @[Mux.scala 31:69:@2561.4]
  wire [15:0] _T_5109; // @[Mux.scala 31:69:@2562.4]
  wire [15:0] _T_5110; // @[Mux.scala 31:69:@2563.4]
  wire [15:0] _T_5111; // @[Mux.scala 31:69:@2564.4]
  wire [15:0] _T_5112; // @[Mux.scala 31:69:@2565.4]
  wire [15:0] _T_5113; // @[Mux.scala 31:69:@2566.4]
  wire [15:0] _T_5114; // @[Mux.scala 31:69:@2567.4]
  wire [15:0] _T_5115; // @[Mux.scala 31:69:@2568.4]
  wire [15:0] _T_5116; // @[Mux.scala 31:69:@2569.4]
  wire [15:0] _T_5117; // @[Mux.scala 31:69:@2570.4]
  wire [15:0] _T_5118; // @[Mux.scala 31:69:@2571.4]
  wire [15:0] _T_5119; // @[Mux.scala 31:69:@2572.4]
  wire [15:0] _T_5120; // @[Mux.scala 31:69:@2573.4]
  wire  _T_5121; // @[OneHot.scala 66:30:@2574.4]
  wire  _T_5122; // @[OneHot.scala 66:30:@2575.4]
  wire  _T_5123; // @[OneHot.scala 66:30:@2576.4]
  wire  _T_5124; // @[OneHot.scala 66:30:@2577.4]
  wire  _T_5125; // @[OneHot.scala 66:30:@2578.4]
  wire  _T_5126; // @[OneHot.scala 66:30:@2579.4]
  wire  _T_5127; // @[OneHot.scala 66:30:@2580.4]
  wire  _T_5128; // @[OneHot.scala 66:30:@2581.4]
  wire  _T_5129; // @[OneHot.scala 66:30:@2582.4]
  wire  _T_5130; // @[OneHot.scala 66:30:@2583.4]
  wire  _T_5131; // @[OneHot.scala 66:30:@2584.4]
  wire  _T_5132; // @[OneHot.scala 66:30:@2585.4]
  wire  _T_5133; // @[OneHot.scala 66:30:@2586.4]
  wire  _T_5134; // @[OneHot.scala 66:30:@2587.4]
  wire  _T_5135; // @[OneHot.scala 66:30:@2588.4]
  wire  _T_5136; // @[OneHot.scala 66:30:@2589.4]
  wire [15:0] _T_5177; // @[Mux.scala 31:69:@2607.4]
  wire [15:0] _T_5178; // @[Mux.scala 31:69:@2608.4]
  wire [15:0] _T_5179; // @[Mux.scala 31:69:@2609.4]
  wire [15:0] _T_5180; // @[Mux.scala 31:69:@2610.4]
  wire [15:0] _T_5181; // @[Mux.scala 31:69:@2611.4]
  wire [15:0] _T_5182; // @[Mux.scala 31:69:@2612.4]
  wire [15:0] _T_5183; // @[Mux.scala 31:69:@2613.4]
  wire [15:0] _T_5184; // @[Mux.scala 31:69:@2614.4]
  wire [15:0] _T_5185; // @[Mux.scala 31:69:@2615.4]
  wire [15:0] _T_5186; // @[Mux.scala 31:69:@2616.4]
  wire [15:0] _T_5187; // @[Mux.scala 31:69:@2617.4]
  wire [15:0] _T_5188; // @[Mux.scala 31:69:@2618.4]
  wire [15:0] _T_5189; // @[Mux.scala 31:69:@2619.4]
  wire [15:0] _T_5190; // @[Mux.scala 31:69:@2620.4]
  wire [15:0] _T_5191; // @[Mux.scala 31:69:@2621.4]
  wire [15:0] _T_5192; // @[Mux.scala 31:69:@2622.4]
  wire  _T_5193; // @[OneHot.scala 66:30:@2623.4]
  wire  _T_5194; // @[OneHot.scala 66:30:@2624.4]
  wire  _T_5195; // @[OneHot.scala 66:30:@2625.4]
  wire  _T_5196; // @[OneHot.scala 66:30:@2626.4]
  wire  _T_5197; // @[OneHot.scala 66:30:@2627.4]
  wire  _T_5198; // @[OneHot.scala 66:30:@2628.4]
  wire  _T_5199; // @[OneHot.scala 66:30:@2629.4]
  wire  _T_5200; // @[OneHot.scala 66:30:@2630.4]
  wire  _T_5201; // @[OneHot.scala 66:30:@2631.4]
  wire  _T_5202; // @[OneHot.scala 66:30:@2632.4]
  wire  _T_5203; // @[OneHot.scala 66:30:@2633.4]
  wire  _T_5204; // @[OneHot.scala 66:30:@2634.4]
  wire  _T_5205; // @[OneHot.scala 66:30:@2635.4]
  wire  _T_5206; // @[OneHot.scala 66:30:@2636.4]
  wire  _T_5207; // @[OneHot.scala 66:30:@2637.4]
  wire  _T_5208; // @[OneHot.scala 66:30:@2638.4]
  wire [15:0] _T_5249; // @[Mux.scala 31:69:@2656.4]
  wire [15:0] _T_5250; // @[Mux.scala 31:69:@2657.4]
  wire [15:0] _T_5251; // @[Mux.scala 31:69:@2658.4]
  wire [15:0] _T_5252; // @[Mux.scala 31:69:@2659.4]
  wire [15:0] _T_5253; // @[Mux.scala 31:69:@2660.4]
  wire [15:0] _T_5254; // @[Mux.scala 31:69:@2661.4]
  wire [15:0] _T_5255; // @[Mux.scala 31:69:@2662.4]
  wire [15:0] _T_5256; // @[Mux.scala 31:69:@2663.4]
  wire [15:0] _T_5257; // @[Mux.scala 31:69:@2664.4]
  wire [15:0] _T_5258; // @[Mux.scala 31:69:@2665.4]
  wire [15:0] _T_5259; // @[Mux.scala 31:69:@2666.4]
  wire [15:0] _T_5260; // @[Mux.scala 31:69:@2667.4]
  wire [15:0] _T_5261; // @[Mux.scala 31:69:@2668.4]
  wire [15:0] _T_5262; // @[Mux.scala 31:69:@2669.4]
  wire [15:0] _T_5263; // @[Mux.scala 31:69:@2670.4]
  wire [15:0] _T_5264; // @[Mux.scala 31:69:@2671.4]
  wire  _T_5265; // @[OneHot.scala 66:30:@2672.4]
  wire  _T_5266; // @[OneHot.scala 66:30:@2673.4]
  wire  _T_5267; // @[OneHot.scala 66:30:@2674.4]
  wire  _T_5268; // @[OneHot.scala 66:30:@2675.4]
  wire  _T_5269; // @[OneHot.scala 66:30:@2676.4]
  wire  _T_5270; // @[OneHot.scala 66:30:@2677.4]
  wire  _T_5271; // @[OneHot.scala 66:30:@2678.4]
  wire  _T_5272; // @[OneHot.scala 66:30:@2679.4]
  wire  _T_5273; // @[OneHot.scala 66:30:@2680.4]
  wire  _T_5274; // @[OneHot.scala 66:30:@2681.4]
  wire  _T_5275; // @[OneHot.scala 66:30:@2682.4]
  wire  _T_5276; // @[OneHot.scala 66:30:@2683.4]
  wire  _T_5277; // @[OneHot.scala 66:30:@2684.4]
  wire  _T_5278; // @[OneHot.scala 66:30:@2685.4]
  wire  _T_5279; // @[OneHot.scala 66:30:@2686.4]
  wire  _T_5280; // @[OneHot.scala 66:30:@2687.4]
  wire [15:0] _T_5321; // @[Mux.scala 31:69:@2705.4]
  wire [15:0] _T_5322; // @[Mux.scala 31:69:@2706.4]
  wire [15:0] _T_5323; // @[Mux.scala 31:69:@2707.4]
  wire [15:0] _T_5324; // @[Mux.scala 31:69:@2708.4]
  wire [15:0] _T_5325; // @[Mux.scala 31:69:@2709.4]
  wire [15:0] _T_5326; // @[Mux.scala 31:69:@2710.4]
  wire [15:0] _T_5327; // @[Mux.scala 31:69:@2711.4]
  wire [15:0] _T_5328; // @[Mux.scala 31:69:@2712.4]
  wire [15:0] _T_5329; // @[Mux.scala 31:69:@2713.4]
  wire [15:0] _T_5330; // @[Mux.scala 31:69:@2714.4]
  wire [15:0] _T_5331; // @[Mux.scala 31:69:@2715.4]
  wire [15:0] _T_5332; // @[Mux.scala 31:69:@2716.4]
  wire [15:0] _T_5333; // @[Mux.scala 31:69:@2717.4]
  wire [15:0] _T_5334; // @[Mux.scala 31:69:@2718.4]
  wire [15:0] _T_5335; // @[Mux.scala 31:69:@2719.4]
  wire [15:0] _T_5336; // @[Mux.scala 31:69:@2720.4]
  wire  _T_5337; // @[OneHot.scala 66:30:@2721.4]
  wire  _T_5338; // @[OneHot.scala 66:30:@2722.4]
  wire  _T_5339; // @[OneHot.scala 66:30:@2723.4]
  wire  _T_5340; // @[OneHot.scala 66:30:@2724.4]
  wire  _T_5341; // @[OneHot.scala 66:30:@2725.4]
  wire  _T_5342; // @[OneHot.scala 66:30:@2726.4]
  wire  _T_5343; // @[OneHot.scala 66:30:@2727.4]
  wire  _T_5344; // @[OneHot.scala 66:30:@2728.4]
  wire  _T_5345; // @[OneHot.scala 66:30:@2729.4]
  wire  _T_5346; // @[OneHot.scala 66:30:@2730.4]
  wire  _T_5347; // @[OneHot.scala 66:30:@2731.4]
  wire  _T_5348; // @[OneHot.scala 66:30:@2732.4]
  wire  _T_5349; // @[OneHot.scala 66:30:@2733.4]
  wire  _T_5350; // @[OneHot.scala 66:30:@2734.4]
  wire  _T_5351; // @[OneHot.scala 66:30:@2735.4]
  wire  _T_5352; // @[OneHot.scala 66:30:@2736.4]
  wire [15:0] _T_5393; // @[Mux.scala 31:69:@2754.4]
  wire [15:0] _T_5394; // @[Mux.scala 31:69:@2755.4]
  wire [15:0] _T_5395; // @[Mux.scala 31:69:@2756.4]
  wire [15:0] _T_5396; // @[Mux.scala 31:69:@2757.4]
  wire [15:0] _T_5397; // @[Mux.scala 31:69:@2758.4]
  wire [15:0] _T_5398; // @[Mux.scala 31:69:@2759.4]
  wire [15:0] _T_5399; // @[Mux.scala 31:69:@2760.4]
  wire [15:0] _T_5400; // @[Mux.scala 31:69:@2761.4]
  wire [15:0] _T_5401; // @[Mux.scala 31:69:@2762.4]
  wire [15:0] _T_5402; // @[Mux.scala 31:69:@2763.4]
  wire [15:0] _T_5403; // @[Mux.scala 31:69:@2764.4]
  wire [15:0] _T_5404; // @[Mux.scala 31:69:@2765.4]
  wire [15:0] _T_5405; // @[Mux.scala 31:69:@2766.4]
  wire [15:0] _T_5406; // @[Mux.scala 31:69:@2767.4]
  wire [15:0] _T_5407; // @[Mux.scala 31:69:@2768.4]
  wire [15:0] _T_5408; // @[Mux.scala 31:69:@2769.4]
  wire  _T_5409; // @[OneHot.scala 66:30:@2770.4]
  wire  _T_5410; // @[OneHot.scala 66:30:@2771.4]
  wire  _T_5411; // @[OneHot.scala 66:30:@2772.4]
  wire  _T_5412; // @[OneHot.scala 66:30:@2773.4]
  wire  _T_5413; // @[OneHot.scala 66:30:@2774.4]
  wire  _T_5414; // @[OneHot.scala 66:30:@2775.4]
  wire  _T_5415; // @[OneHot.scala 66:30:@2776.4]
  wire  _T_5416; // @[OneHot.scala 66:30:@2777.4]
  wire  _T_5417; // @[OneHot.scala 66:30:@2778.4]
  wire  _T_5418; // @[OneHot.scala 66:30:@2779.4]
  wire  _T_5419; // @[OneHot.scala 66:30:@2780.4]
  wire  _T_5420; // @[OneHot.scala 66:30:@2781.4]
  wire  _T_5421; // @[OneHot.scala 66:30:@2782.4]
  wire  _T_5422; // @[OneHot.scala 66:30:@2783.4]
  wire  _T_5423; // @[OneHot.scala 66:30:@2784.4]
  wire  _T_5424; // @[OneHot.scala 66:30:@2785.4]
  wire [7:0] _T_5489; // @[Mux.scala 19:72:@2809.4]
  wire [15:0] _T_5497; // @[Mux.scala 19:72:@2817.4]
  wire [15:0] _T_5499; // @[Mux.scala 19:72:@2818.4]
  wire [7:0] _T_5506; // @[Mux.scala 19:72:@2825.4]
  wire [15:0] _T_5514; // @[Mux.scala 19:72:@2833.4]
  wire [15:0] _T_5516; // @[Mux.scala 19:72:@2834.4]
  wire [7:0] _T_5523; // @[Mux.scala 19:72:@2841.4]
  wire [15:0] _T_5531; // @[Mux.scala 19:72:@2849.4]
  wire [15:0] _T_5533; // @[Mux.scala 19:72:@2850.4]
  wire [7:0] _T_5540; // @[Mux.scala 19:72:@2857.4]
  wire [15:0] _T_5548; // @[Mux.scala 19:72:@2865.4]
  wire [15:0] _T_5550; // @[Mux.scala 19:72:@2866.4]
  wire [7:0] _T_5557; // @[Mux.scala 19:72:@2873.4]
  wire [15:0] _T_5565; // @[Mux.scala 19:72:@2881.4]
  wire [15:0] _T_5567; // @[Mux.scala 19:72:@2882.4]
  wire [7:0] _T_5574; // @[Mux.scala 19:72:@2889.4]
  wire [15:0] _T_5582; // @[Mux.scala 19:72:@2897.4]
  wire [15:0] _T_5584; // @[Mux.scala 19:72:@2898.4]
  wire [7:0] _T_5591; // @[Mux.scala 19:72:@2905.4]
  wire [15:0] _T_5599; // @[Mux.scala 19:72:@2913.4]
  wire [15:0] _T_5601; // @[Mux.scala 19:72:@2914.4]
  wire [7:0] _T_5608; // @[Mux.scala 19:72:@2921.4]
  wire [15:0] _T_5616; // @[Mux.scala 19:72:@2929.4]
  wire [15:0] _T_5618; // @[Mux.scala 19:72:@2930.4]
  wire [7:0] _T_5625; // @[Mux.scala 19:72:@2937.4]
  wire [15:0] _T_5633; // @[Mux.scala 19:72:@2945.4]
  wire [15:0] _T_5635; // @[Mux.scala 19:72:@2946.4]
  wire [7:0] _T_5642; // @[Mux.scala 19:72:@2953.4]
  wire [15:0] _T_5650; // @[Mux.scala 19:72:@2961.4]
  wire [15:0] _T_5652; // @[Mux.scala 19:72:@2962.4]
  wire [7:0] _T_5659; // @[Mux.scala 19:72:@2969.4]
  wire [15:0] _T_5667; // @[Mux.scala 19:72:@2977.4]
  wire [15:0] _T_5669; // @[Mux.scala 19:72:@2978.4]
  wire [7:0] _T_5676; // @[Mux.scala 19:72:@2985.4]
  wire [15:0] _T_5684; // @[Mux.scala 19:72:@2993.4]
  wire [15:0] _T_5686; // @[Mux.scala 19:72:@2994.4]
  wire [7:0] _T_5693; // @[Mux.scala 19:72:@3001.4]
  wire [15:0] _T_5701; // @[Mux.scala 19:72:@3009.4]
  wire [15:0] _T_5703; // @[Mux.scala 19:72:@3010.4]
  wire [7:0] _T_5710; // @[Mux.scala 19:72:@3017.4]
  wire [15:0] _T_5718; // @[Mux.scala 19:72:@3025.4]
  wire [15:0] _T_5720; // @[Mux.scala 19:72:@3026.4]
  wire [7:0] _T_5727; // @[Mux.scala 19:72:@3033.4]
  wire [15:0] _T_5735; // @[Mux.scala 19:72:@3041.4]
  wire [15:0] _T_5737; // @[Mux.scala 19:72:@3042.4]
  wire [7:0] _T_5744; // @[Mux.scala 19:72:@3049.4]
  wire [15:0] _T_5752; // @[Mux.scala 19:72:@3057.4]
  wire [15:0] _T_5754; // @[Mux.scala 19:72:@3058.4]
  wire [15:0] _T_5755; // @[Mux.scala 19:72:@3059.4]
  wire [15:0] _T_5756; // @[Mux.scala 19:72:@3060.4]
  wire [15:0] _T_5757; // @[Mux.scala 19:72:@3061.4]
  wire [15:0] _T_5758; // @[Mux.scala 19:72:@3062.4]
  wire [15:0] _T_5759; // @[Mux.scala 19:72:@3063.4]
  wire [15:0] _T_5760; // @[Mux.scala 19:72:@3064.4]
  wire [15:0] _T_5761; // @[Mux.scala 19:72:@3065.4]
  wire [15:0] _T_5762; // @[Mux.scala 19:72:@3066.4]
  wire [15:0] _T_5763; // @[Mux.scala 19:72:@3067.4]
  wire [15:0] _T_5764; // @[Mux.scala 19:72:@3068.4]
  wire [15:0] _T_5765; // @[Mux.scala 19:72:@3069.4]
  wire [15:0] _T_5766; // @[Mux.scala 19:72:@3070.4]
  wire [15:0] _T_5767; // @[Mux.scala 19:72:@3071.4]
  wire [15:0] _T_5768; // @[Mux.scala 19:72:@3072.4]
  wire [15:0] _T_5769; // @[Mux.scala 19:72:@3073.4]
  wire  inputAddrPriorityPorts_0_0; // @[Mux.scala 19:72:@3077.4]
  wire  inputAddrPriorityPorts_0_1; // @[Mux.scala 19:72:@3079.4]
  wire  inputAddrPriorityPorts_0_2; // @[Mux.scala 19:72:@3081.4]
  wire  inputAddrPriorityPorts_0_3; // @[Mux.scala 19:72:@3083.4]
  wire  inputAddrPriorityPorts_0_4; // @[Mux.scala 19:72:@3085.4]
  wire  inputAddrPriorityPorts_0_5; // @[Mux.scala 19:72:@3087.4]
  wire  inputAddrPriorityPorts_0_6; // @[Mux.scala 19:72:@3089.4]
  wire  inputAddrPriorityPorts_0_7; // @[Mux.scala 19:72:@3091.4]
  wire  inputAddrPriorityPorts_0_8; // @[Mux.scala 19:72:@3093.4]
  wire  inputAddrPriorityPorts_0_9; // @[Mux.scala 19:72:@3095.4]
  wire  inputAddrPriorityPorts_0_10; // @[Mux.scala 19:72:@3097.4]
  wire  inputAddrPriorityPorts_0_11; // @[Mux.scala 19:72:@3099.4]
  wire  inputAddrPriorityPorts_0_12; // @[Mux.scala 19:72:@3101.4]
  wire  inputAddrPriorityPorts_0_13; // @[Mux.scala 19:72:@3103.4]
  wire  inputAddrPriorityPorts_0_14; // @[Mux.scala 19:72:@3105.4]
  wire  inputAddrPriorityPorts_0_15; // @[Mux.scala 19:72:@3107.4]
  wire [15:0] _T_5971; // @[Mux.scala 31:69:@3161.4]
  wire [15:0] _T_5972; // @[Mux.scala 31:69:@3162.4]
  wire [15:0] _T_5973; // @[Mux.scala 31:69:@3163.4]
  wire [15:0] _T_5974; // @[Mux.scala 31:69:@3164.4]
  wire [15:0] _T_5975; // @[Mux.scala 31:69:@3165.4]
  wire [15:0] _T_5976; // @[Mux.scala 31:69:@3166.4]
  wire [15:0] _T_5977; // @[Mux.scala 31:69:@3167.4]
  wire [15:0] _T_5978; // @[Mux.scala 31:69:@3168.4]
  wire [15:0] _T_5979; // @[Mux.scala 31:69:@3169.4]
  wire [15:0] _T_5980; // @[Mux.scala 31:69:@3170.4]
  wire [15:0] _T_5981; // @[Mux.scala 31:69:@3171.4]
  wire [15:0] _T_5982; // @[Mux.scala 31:69:@3172.4]
  wire [15:0] _T_5983; // @[Mux.scala 31:69:@3173.4]
  wire [15:0] _T_5984; // @[Mux.scala 31:69:@3174.4]
  wire [15:0] _T_5985; // @[Mux.scala 31:69:@3175.4]
  wire [15:0] _T_5986; // @[Mux.scala 31:69:@3176.4]
  wire  _T_5987; // @[OneHot.scala 66:30:@3177.4]
  wire  _T_5988; // @[OneHot.scala 66:30:@3178.4]
  wire  _T_5989; // @[OneHot.scala 66:30:@3179.4]
  wire  _T_5990; // @[OneHot.scala 66:30:@3180.4]
  wire  _T_5991; // @[OneHot.scala 66:30:@3181.4]
  wire  _T_5992; // @[OneHot.scala 66:30:@3182.4]
  wire  _T_5993; // @[OneHot.scala 66:30:@3183.4]
  wire  _T_5994; // @[OneHot.scala 66:30:@3184.4]
  wire  _T_5995; // @[OneHot.scala 66:30:@3185.4]
  wire  _T_5996; // @[OneHot.scala 66:30:@3186.4]
  wire  _T_5997; // @[OneHot.scala 66:30:@3187.4]
  wire  _T_5998; // @[OneHot.scala 66:30:@3188.4]
  wire  _T_5999; // @[OneHot.scala 66:30:@3189.4]
  wire  _T_6000; // @[OneHot.scala 66:30:@3190.4]
  wire  _T_6001; // @[OneHot.scala 66:30:@3191.4]
  wire  _T_6002; // @[OneHot.scala 66:30:@3192.4]
  wire [15:0] _T_6043; // @[Mux.scala 31:69:@3210.4]
  wire [15:0] _T_6044; // @[Mux.scala 31:69:@3211.4]
  wire [15:0] _T_6045; // @[Mux.scala 31:69:@3212.4]
  wire [15:0] _T_6046; // @[Mux.scala 31:69:@3213.4]
  wire [15:0] _T_6047; // @[Mux.scala 31:69:@3214.4]
  wire [15:0] _T_6048; // @[Mux.scala 31:69:@3215.4]
  wire [15:0] _T_6049; // @[Mux.scala 31:69:@3216.4]
  wire [15:0] _T_6050; // @[Mux.scala 31:69:@3217.4]
  wire [15:0] _T_6051; // @[Mux.scala 31:69:@3218.4]
  wire [15:0] _T_6052; // @[Mux.scala 31:69:@3219.4]
  wire [15:0] _T_6053; // @[Mux.scala 31:69:@3220.4]
  wire [15:0] _T_6054; // @[Mux.scala 31:69:@3221.4]
  wire [15:0] _T_6055; // @[Mux.scala 31:69:@3222.4]
  wire [15:0] _T_6056; // @[Mux.scala 31:69:@3223.4]
  wire [15:0] _T_6057; // @[Mux.scala 31:69:@3224.4]
  wire [15:0] _T_6058; // @[Mux.scala 31:69:@3225.4]
  wire  _T_6059; // @[OneHot.scala 66:30:@3226.4]
  wire  _T_6060; // @[OneHot.scala 66:30:@3227.4]
  wire  _T_6061; // @[OneHot.scala 66:30:@3228.4]
  wire  _T_6062; // @[OneHot.scala 66:30:@3229.4]
  wire  _T_6063; // @[OneHot.scala 66:30:@3230.4]
  wire  _T_6064; // @[OneHot.scala 66:30:@3231.4]
  wire  _T_6065; // @[OneHot.scala 66:30:@3232.4]
  wire  _T_6066; // @[OneHot.scala 66:30:@3233.4]
  wire  _T_6067; // @[OneHot.scala 66:30:@3234.4]
  wire  _T_6068; // @[OneHot.scala 66:30:@3235.4]
  wire  _T_6069; // @[OneHot.scala 66:30:@3236.4]
  wire  _T_6070; // @[OneHot.scala 66:30:@3237.4]
  wire  _T_6071; // @[OneHot.scala 66:30:@3238.4]
  wire  _T_6072; // @[OneHot.scala 66:30:@3239.4]
  wire  _T_6073; // @[OneHot.scala 66:30:@3240.4]
  wire  _T_6074; // @[OneHot.scala 66:30:@3241.4]
  wire [15:0] _T_6115; // @[Mux.scala 31:69:@3259.4]
  wire [15:0] _T_6116; // @[Mux.scala 31:69:@3260.4]
  wire [15:0] _T_6117; // @[Mux.scala 31:69:@3261.4]
  wire [15:0] _T_6118; // @[Mux.scala 31:69:@3262.4]
  wire [15:0] _T_6119; // @[Mux.scala 31:69:@3263.4]
  wire [15:0] _T_6120; // @[Mux.scala 31:69:@3264.4]
  wire [15:0] _T_6121; // @[Mux.scala 31:69:@3265.4]
  wire [15:0] _T_6122; // @[Mux.scala 31:69:@3266.4]
  wire [15:0] _T_6123; // @[Mux.scala 31:69:@3267.4]
  wire [15:0] _T_6124; // @[Mux.scala 31:69:@3268.4]
  wire [15:0] _T_6125; // @[Mux.scala 31:69:@3269.4]
  wire [15:0] _T_6126; // @[Mux.scala 31:69:@3270.4]
  wire [15:0] _T_6127; // @[Mux.scala 31:69:@3271.4]
  wire [15:0] _T_6128; // @[Mux.scala 31:69:@3272.4]
  wire [15:0] _T_6129; // @[Mux.scala 31:69:@3273.4]
  wire [15:0] _T_6130; // @[Mux.scala 31:69:@3274.4]
  wire  _T_6131; // @[OneHot.scala 66:30:@3275.4]
  wire  _T_6132; // @[OneHot.scala 66:30:@3276.4]
  wire  _T_6133; // @[OneHot.scala 66:30:@3277.4]
  wire  _T_6134; // @[OneHot.scala 66:30:@3278.4]
  wire  _T_6135; // @[OneHot.scala 66:30:@3279.4]
  wire  _T_6136; // @[OneHot.scala 66:30:@3280.4]
  wire  _T_6137; // @[OneHot.scala 66:30:@3281.4]
  wire  _T_6138; // @[OneHot.scala 66:30:@3282.4]
  wire  _T_6139; // @[OneHot.scala 66:30:@3283.4]
  wire  _T_6140; // @[OneHot.scala 66:30:@3284.4]
  wire  _T_6141; // @[OneHot.scala 66:30:@3285.4]
  wire  _T_6142; // @[OneHot.scala 66:30:@3286.4]
  wire  _T_6143; // @[OneHot.scala 66:30:@3287.4]
  wire  _T_6144; // @[OneHot.scala 66:30:@3288.4]
  wire  _T_6145; // @[OneHot.scala 66:30:@3289.4]
  wire  _T_6146; // @[OneHot.scala 66:30:@3290.4]
  wire [15:0] _T_6187; // @[Mux.scala 31:69:@3308.4]
  wire [15:0] _T_6188; // @[Mux.scala 31:69:@3309.4]
  wire [15:0] _T_6189; // @[Mux.scala 31:69:@3310.4]
  wire [15:0] _T_6190; // @[Mux.scala 31:69:@3311.4]
  wire [15:0] _T_6191; // @[Mux.scala 31:69:@3312.4]
  wire [15:0] _T_6192; // @[Mux.scala 31:69:@3313.4]
  wire [15:0] _T_6193; // @[Mux.scala 31:69:@3314.4]
  wire [15:0] _T_6194; // @[Mux.scala 31:69:@3315.4]
  wire [15:0] _T_6195; // @[Mux.scala 31:69:@3316.4]
  wire [15:0] _T_6196; // @[Mux.scala 31:69:@3317.4]
  wire [15:0] _T_6197; // @[Mux.scala 31:69:@3318.4]
  wire [15:0] _T_6198; // @[Mux.scala 31:69:@3319.4]
  wire [15:0] _T_6199; // @[Mux.scala 31:69:@3320.4]
  wire [15:0] _T_6200; // @[Mux.scala 31:69:@3321.4]
  wire [15:0] _T_6201; // @[Mux.scala 31:69:@3322.4]
  wire [15:0] _T_6202; // @[Mux.scala 31:69:@3323.4]
  wire  _T_6203; // @[OneHot.scala 66:30:@3324.4]
  wire  _T_6204; // @[OneHot.scala 66:30:@3325.4]
  wire  _T_6205; // @[OneHot.scala 66:30:@3326.4]
  wire  _T_6206; // @[OneHot.scala 66:30:@3327.4]
  wire  _T_6207; // @[OneHot.scala 66:30:@3328.4]
  wire  _T_6208; // @[OneHot.scala 66:30:@3329.4]
  wire  _T_6209; // @[OneHot.scala 66:30:@3330.4]
  wire  _T_6210; // @[OneHot.scala 66:30:@3331.4]
  wire  _T_6211; // @[OneHot.scala 66:30:@3332.4]
  wire  _T_6212; // @[OneHot.scala 66:30:@3333.4]
  wire  _T_6213; // @[OneHot.scala 66:30:@3334.4]
  wire  _T_6214; // @[OneHot.scala 66:30:@3335.4]
  wire  _T_6215; // @[OneHot.scala 66:30:@3336.4]
  wire  _T_6216; // @[OneHot.scala 66:30:@3337.4]
  wire  _T_6217; // @[OneHot.scala 66:30:@3338.4]
  wire  _T_6218; // @[OneHot.scala 66:30:@3339.4]
  wire [15:0] _T_6259; // @[Mux.scala 31:69:@3357.4]
  wire [15:0] _T_6260; // @[Mux.scala 31:69:@3358.4]
  wire [15:0] _T_6261; // @[Mux.scala 31:69:@3359.4]
  wire [15:0] _T_6262; // @[Mux.scala 31:69:@3360.4]
  wire [15:0] _T_6263; // @[Mux.scala 31:69:@3361.4]
  wire [15:0] _T_6264; // @[Mux.scala 31:69:@3362.4]
  wire [15:0] _T_6265; // @[Mux.scala 31:69:@3363.4]
  wire [15:0] _T_6266; // @[Mux.scala 31:69:@3364.4]
  wire [15:0] _T_6267; // @[Mux.scala 31:69:@3365.4]
  wire [15:0] _T_6268; // @[Mux.scala 31:69:@3366.4]
  wire [15:0] _T_6269; // @[Mux.scala 31:69:@3367.4]
  wire [15:0] _T_6270; // @[Mux.scala 31:69:@3368.4]
  wire [15:0] _T_6271; // @[Mux.scala 31:69:@3369.4]
  wire [15:0] _T_6272; // @[Mux.scala 31:69:@3370.4]
  wire [15:0] _T_6273; // @[Mux.scala 31:69:@3371.4]
  wire [15:0] _T_6274; // @[Mux.scala 31:69:@3372.4]
  wire  _T_6275; // @[OneHot.scala 66:30:@3373.4]
  wire  _T_6276; // @[OneHot.scala 66:30:@3374.4]
  wire  _T_6277; // @[OneHot.scala 66:30:@3375.4]
  wire  _T_6278; // @[OneHot.scala 66:30:@3376.4]
  wire  _T_6279; // @[OneHot.scala 66:30:@3377.4]
  wire  _T_6280; // @[OneHot.scala 66:30:@3378.4]
  wire  _T_6281; // @[OneHot.scala 66:30:@3379.4]
  wire  _T_6282; // @[OneHot.scala 66:30:@3380.4]
  wire  _T_6283; // @[OneHot.scala 66:30:@3381.4]
  wire  _T_6284; // @[OneHot.scala 66:30:@3382.4]
  wire  _T_6285; // @[OneHot.scala 66:30:@3383.4]
  wire  _T_6286; // @[OneHot.scala 66:30:@3384.4]
  wire  _T_6287; // @[OneHot.scala 66:30:@3385.4]
  wire  _T_6288; // @[OneHot.scala 66:30:@3386.4]
  wire  _T_6289; // @[OneHot.scala 66:30:@3387.4]
  wire  _T_6290; // @[OneHot.scala 66:30:@3388.4]
  wire [15:0] _T_6331; // @[Mux.scala 31:69:@3406.4]
  wire [15:0] _T_6332; // @[Mux.scala 31:69:@3407.4]
  wire [15:0] _T_6333; // @[Mux.scala 31:69:@3408.4]
  wire [15:0] _T_6334; // @[Mux.scala 31:69:@3409.4]
  wire [15:0] _T_6335; // @[Mux.scala 31:69:@3410.4]
  wire [15:0] _T_6336; // @[Mux.scala 31:69:@3411.4]
  wire [15:0] _T_6337; // @[Mux.scala 31:69:@3412.4]
  wire [15:0] _T_6338; // @[Mux.scala 31:69:@3413.4]
  wire [15:0] _T_6339; // @[Mux.scala 31:69:@3414.4]
  wire [15:0] _T_6340; // @[Mux.scala 31:69:@3415.4]
  wire [15:0] _T_6341; // @[Mux.scala 31:69:@3416.4]
  wire [15:0] _T_6342; // @[Mux.scala 31:69:@3417.4]
  wire [15:0] _T_6343; // @[Mux.scala 31:69:@3418.4]
  wire [15:0] _T_6344; // @[Mux.scala 31:69:@3419.4]
  wire [15:0] _T_6345; // @[Mux.scala 31:69:@3420.4]
  wire [15:0] _T_6346; // @[Mux.scala 31:69:@3421.4]
  wire  _T_6347; // @[OneHot.scala 66:30:@3422.4]
  wire  _T_6348; // @[OneHot.scala 66:30:@3423.4]
  wire  _T_6349; // @[OneHot.scala 66:30:@3424.4]
  wire  _T_6350; // @[OneHot.scala 66:30:@3425.4]
  wire  _T_6351; // @[OneHot.scala 66:30:@3426.4]
  wire  _T_6352; // @[OneHot.scala 66:30:@3427.4]
  wire  _T_6353; // @[OneHot.scala 66:30:@3428.4]
  wire  _T_6354; // @[OneHot.scala 66:30:@3429.4]
  wire  _T_6355; // @[OneHot.scala 66:30:@3430.4]
  wire  _T_6356; // @[OneHot.scala 66:30:@3431.4]
  wire  _T_6357; // @[OneHot.scala 66:30:@3432.4]
  wire  _T_6358; // @[OneHot.scala 66:30:@3433.4]
  wire  _T_6359; // @[OneHot.scala 66:30:@3434.4]
  wire  _T_6360; // @[OneHot.scala 66:30:@3435.4]
  wire  _T_6361; // @[OneHot.scala 66:30:@3436.4]
  wire  _T_6362; // @[OneHot.scala 66:30:@3437.4]
  wire [15:0] _T_6403; // @[Mux.scala 31:69:@3455.4]
  wire [15:0] _T_6404; // @[Mux.scala 31:69:@3456.4]
  wire [15:0] _T_6405; // @[Mux.scala 31:69:@3457.4]
  wire [15:0] _T_6406; // @[Mux.scala 31:69:@3458.4]
  wire [15:0] _T_6407; // @[Mux.scala 31:69:@3459.4]
  wire [15:0] _T_6408; // @[Mux.scala 31:69:@3460.4]
  wire [15:0] _T_6409; // @[Mux.scala 31:69:@3461.4]
  wire [15:0] _T_6410; // @[Mux.scala 31:69:@3462.4]
  wire [15:0] _T_6411; // @[Mux.scala 31:69:@3463.4]
  wire [15:0] _T_6412; // @[Mux.scala 31:69:@3464.4]
  wire [15:0] _T_6413; // @[Mux.scala 31:69:@3465.4]
  wire [15:0] _T_6414; // @[Mux.scala 31:69:@3466.4]
  wire [15:0] _T_6415; // @[Mux.scala 31:69:@3467.4]
  wire [15:0] _T_6416; // @[Mux.scala 31:69:@3468.4]
  wire [15:0] _T_6417; // @[Mux.scala 31:69:@3469.4]
  wire [15:0] _T_6418; // @[Mux.scala 31:69:@3470.4]
  wire  _T_6419; // @[OneHot.scala 66:30:@3471.4]
  wire  _T_6420; // @[OneHot.scala 66:30:@3472.4]
  wire  _T_6421; // @[OneHot.scala 66:30:@3473.4]
  wire  _T_6422; // @[OneHot.scala 66:30:@3474.4]
  wire  _T_6423; // @[OneHot.scala 66:30:@3475.4]
  wire  _T_6424; // @[OneHot.scala 66:30:@3476.4]
  wire  _T_6425; // @[OneHot.scala 66:30:@3477.4]
  wire  _T_6426; // @[OneHot.scala 66:30:@3478.4]
  wire  _T_6427; // @[OneHot.scala 66:30:@3479.4]
  wire  _T_6428; // @[OneHot.scala 66:30:@3480.4]
  wire  _T_6429; // @[OneHot.scala 66:30:@3481.4]
  wire  _T_6430; // @[OneHot.scala 66:30:@3482.4]
  wire  _T_6431; // @[OneHot.scala 66:30:@3483.4]
  wire  _T_6432; // @[OneHot.scala 66:30:@3484.4]
  wire  _T_6433; // @[OneHot.scala 66:30:@3485.4]
  wire  _T_6434; // @[OneHot.scala 66:30:@3486.4]
  wire [15:0] _T_6475; // @[Mux.scala 31:69:@3504.4]
  wire [15:0] _T_6476; // @[Mux.scala 31:69:@3505.4]
  wire [15:0] _T_6477; // @[Mux.scala 31:69:@3506.4]
  wire [15:0] _T_6478; // @[Mux.scala 31:69:@3507.4]
  wire [15:0] _T_6479; // @[Mux.scala 31:69:@3508.4]
  wire [15:0] _T_6480; // @[Mux.scala 31:69:@3509.4]
  wire [15:0] _T_6481; // @[Mux.scala 31:69:@3510.4]
  wire [15:0] _T_6482; // @[Mux.scala 31:69:@3511.4]
  wire [15:0] _T_6483; // @[Mux.scala 31:69:@3512.4]
  wire [15:0] _T_6484; // @[Mux.scala 31:69:@3513.4]
  wire [15:0] _T_6485; // @[Mux.scala 31:69:@3514.4]
  wire [15:0] _T_6486; // @[Mux.scala 31:69:@3515.4]
  wire [15:0] _T_6487; // @[Mux.scala 31:69:@3516.4]
  wire [15:0] _T_6488; // @[Mux.scala 31:69:@3517.4]
  wire [15:0] _T_6489; // @[Mux.scala 31:69:@3518.4]
  wire [15:0] _T_6490; // @[Mux.scala 31:69:@3519.4]
  wire  _T_6491; // @[OneHot.scala 66:30:@3520.4]
  wire  _T_6492; // @[OneHot.scala 66:30:@3521.4]
  wire  _T_6493; // @[OneHot.scala 66:30:@3522.4]
  wire  _T_6494; // @[OneHot.scala 66:30:@3523.4]
  wire  _T_6495; // @[OneHot.scala 66:30:@3524.4]
  wire  _T_6496; // @[OneHot.scala 66:30:@3525.4]
  wire  _T_6497; // @[OneHot.scala 66:30:@3526.4]
  wire  _T_6498; // @[OneHot.scala 66:30:@3527.4]
  wire  _T_6499; // @[OneHot.scala 66:30:@3528.4]
  wire  _T_6500; // @[OneHot.scala 66:30:@3529.4]
  wire  _T_6501; // @[OneHot.scala 66:30:@3530.4]
  wire  _T_6502; // @[OneHot.scala 66:30:@3531.4]
  wire  _T_6503; // @[OneHot.scala 66:30:@3532.4]
  wire  _T_6504; // @[OneHot.scala 66:30:@3533.4]
  wire  _T_6505; // @[OneHot.scala 66:30:@3534.4]
  wire  _T_6506; // @[OneHot.scala 66:30:@3535.4]
  wire [15:0] _T_6547; // @[Mux.scala 31:69:@3553.4]
  wire [15:0] _T_6548; // @[Mux.scala 31:69:@3554.4]
  wire [15:0] _T_6549; // @[Mux.scala 31:69:@3555.4]
  wire [15:0] _T_6550; // @[Mux.scala 31:69:@3556.4]
  wire [15:0] _T_6551; // @[Mux.scala 31:69:@3557.4]
  wire [15:0] _T_6552; // @[Mux.scala 31:69:@3558.4]
  wire [15:0] _T_6553; // @[Mux.scala 31:69:@3559.4]
  wire [15:0] _T_6554; // @[Mux.scala 31:69:@3560.4]
  wire [15:0] _T_6555; // @[Mux.scala 31:69:@3561.4]
  wire [15:0] _T_6556; // @[Mux.scala 31:69:@3562.4]
  wire [15:0] _T_6557; // @[Mux.scala 31:69:@3563.4]
  wire [15:0] _T_6558; // @[Mux.scala 31:69:@3564.4]
  wire [15:0] _T_6559; // @[Mux.scala 31:69:@3565.4]
  wire [15:0] _T_6560; // @[Mux.scala 31:69:@3566.4]
  wire [15:0] _T_6561; // @[Mux.scala 31:69:@3567.4]
  wire [15:0] _T_6562; // @[Mux.scala 31:69:@3568.4]
  wire  _T_6563; // @[OneHot.scala 66:30:@3569.4]
  wire  _T_6564; // @[OneHot.scala 66:30:@3570.4]
  wire  _T_6565; // @[OneHot.scala 66:30:@3571.4]
  wire  _T_6566; // @[OneHot.scala 66:30:@3572.4]
  wire  _T_6567; // @[OneHot.scala 66:30:@3573.4]
  wire  _T_6568; // @[OneHot.scala 66:30:@3574.4]
  wire  _T_6569; // @[OneHot.scala 66:30:@3575.4]
  wire  _T_6570; // @[OneHot.scala 66:30:@3576.4]
  wire  _T_6571; // @[OneHot.scala 66:30:@3577.4]
  wire  _T_6572; // @[OneHot.scala 66:30:@3578.4]
  wire  _T_6573; // @[OneHot.scala 66:30:@3579.4]
  wire  _T_6574; // @[OneHot.scala 66:30:@3580.4]
  wire  _T_6575; // @[OneHot.scala 66:30:@3581.4]
  wire  _T_6576; // @[OneHot.scala 66:30:@3582.4]
  wire  _T_6577; // @[OneHot.scala 66:30:@3583.4]
  wire  _T_6578; // @[OneHot.scala 66:30:@3584.4]
  wire [15:0] _T_6619; // @[Mux.scala 31:69:@3602.4]
  wire [15:0] _T_6620; // @[Mux.scala 31:69:@3603.4]
  wire [15:0] _T_6621; // @[Mux.scala 31:69:@3604.4]
  wire [15:0] _T_6622; // @[Mux.scala 31:69:@3605.4]
  wire [15:0] _T_6623; // @[Mux.scala 31:69:@3606.4]
  wire [15:0] _T_6624; // @[Mux.scala 31:69:@3607.4]
  wire [15:0] _T_6625; // @[Mux.scala 31:69:@3608.4]
  wire [15:0] _T_6626; // @[Mux.scala 31:69:@3609.4]
  wire [15:0] _T_6627; // @[Mux.scala 31:69:@3610.4]
  wire [15:0] _T_6628; // @[Mux.scala 31:69:@3611.4]
  wire [15:0] _T_6629; // @[Mux.scala 31:69:@3612.4]
  wire [15:0] _T_6630; // @[Mux.scala 31:69:@3613.4]
  wire [15:0] _T_6631; // @[Mux.scala 31:69:@3614.4]
  wire [15:0] _T_6632; // @[Mux.scala 31:69:@3615.4]
  wire [15:0] _T_6633; // @[Mux.scala 31:69:@3616.4]
  wire [15:0] _T_6634; // @[Mux.scala 31:69:@3617.4]
  wire  _T_6635; // @[OneHot.scala 66:30:@3618.4]
  wire  _T_6636; // @[OneHot.scala 66:30:@3619.4]
  wire  _T_6637; // @[OneHot.scala 66:30:@3620.4]
  wire  _T_6638; // @[OneHot.scala 66:30:@3621.4]
  wire  _T_6639; // @[OneHot.scala 66:30:@3622.4]
  wire  _T_6640; // @[OneHot.scala 66:30:@3623.4]
  wire  _T_6641; // @[OneHot.scala 66:30:@3624.4]
  wire  _T_6642; // @[OneHot.scala 66:30:@3625.4]
  wire  _T_6643; // @[OneHot.scala 66:30:@3626.4]
  wire  _T_6644; // @[OneHot.scala 66:30:@3627.4]
  wire  _T_6645; // @[OneHot.scala 66:30:@3628.4]
  wire  _T_6646; // @[OneHot.scala 66:30:@3629.4]
  wire  _T_6647; // @[OneHot.scala 66:30:@3630.4]
  wire  _T_6648; // @[OneHot.scala 66:30:@3631.4]
  wire  _T_6649; // @[OneHot.scala 66:30:@3632.4]
  wire  _T_6650; // @[OneHot.scala 66:30:@3633.4]
  wire [15:0] _T_6691; // @[Mux.scala 31:69:@3651.4]
  wire [15:0] _T_6692; // @[Mux.scala 31:69:@3652.4]
  wire [15:0] _T_6693; // @[Mux.scala 31:69:@3653.4]
  wire [15:0] _T_6694; // @[Mux.scala 31:69:@3654.4]
  wire [15:0] _T_6695; // @[Mux.scala 31:69:@3655.4]
  wire [15:0] _T_6696; // @[Mux.scala 31:69:@3656.4]
  wire [15:0] _T_6697; // @[Mux.scala 31:69:@3657.4]
  wire [15:0] _T_6698; // @[Mux.scala 31:69:@3658.4]
  wire [15:0] _T_6699; // @[Mux.scala 31:69:@3659.4]
  wire [15:0] _T_6700; // @[Mux.scala 31:69:@3660.4]
  wire [15:0] _T_6701; // @[Mux.scala 31:69:@3661.4]
  wire [15:0] _T_6702; // @[Mux.scala 31:69:@3662.4]
  wire [15:0] _T_6703; // @[Mux.scala 31:69:@3663.4]
  wire [15:0] _T_6704; // @[Mux.scala 31:69:@3664.4]
  wire [15:0] _T_6705; // @[Mux.scala 31:69:@3665.4]
  wire [15:0] _T_6706; // @[Mux.scala 31:69:@3666.4]
  wire  _T_6707; // @[OneHot.scala 66:30:@3667.4]
  wire  _T_6708; // @[OneHot.scala 66:30:@3668.4]
  wire  _T_6709; // @[OneHot.scala 66:30:@3669.4]
  wire  _T_6710; // @[OneHot.scala 66:30:@3670.4]
  wire  _T_6711; // @[OneHot.scala 66:30:@3671.4]
  wire  _T_6712; // @[OneHot.scala 66:30:@3672.4]
  wire  _T_6713; // @[OneHot.scala 66:30:@3673.4]
  wire  _T_6714; // @[OneHot.scala 66:30:@3674.4]
  wire  _T_6715; // @[OneHot.scala 66:30:@3675.4]
  wire  _T_6716; // @[OneHot.scala 66:30:@3676.4]
  wire  _T_6717; // @[OneHot.scala 66:30:@3677.4]
  wire  _T_6718; // @[OneHot.scala 66:30:@3678.4]
  wire  _T_6719; // @[OneHot.scala 66:30:@3679.4]
  wire  _T_6720; // @[OneHot.scala 66:30:@3680.4]
  wire  _T_6721; // @[OneHot.scala 66:30:@3681.4]
  wire  _T_6722; // @[OneHot.scala 66:30:@3682.4]
  wire [15:0] _T_6763; // @[Mux.scala 31:69:@3700.4]
  wire [15:0] _T_6764; // @[Mux.scala 31:69:@3701.4]
  wire [15:0] _T_6765; // @[Mux.scala 31:69:@3702.4]
  wire [15:0] _T_6766; // @[Mux.scala 31:69:@3703.4]
  wire [15:0] _T_6767; // @[Mux.scala 31:69:@3704.4]
  wire [15:0] _T_6768; // @[Mux.scala 31:69:@3705.4]
  wire [15:0] _T_6769; // @[Mux.scala 31:69:@3706.4]
  wire [15:0] _T_6770; // @[Mux.scala 31:69:@3707.4]
  wire [15:0] _T_6771; // @[Mux.scala 31:69:@3708.4]
  wire [15:0] _T_6772; // @[Mux.scala 31:69:@3709.4]
  wire [15:0] _T_6773; // @[Mux.scala 31:69:@3710.4]
  wire [15:0] _T_6774; // @[Mux.scala 31:69:@3711.4]
  wire [15:0] _T_6775; // @[Mux.scala 31:69:@3712.4]
  wire [15:0] _T_6776; // @[Mux.scala 31:69:@3713.4]
  wire [15:0] _T_6777; // @[Mux.scala 31:69:@3714.4]
  wire [15:0] _T_6778; // @[Mux.scala 31:69:@3715.4]
  wire  _T_6779; // @[OneHot.scala 66:30:@3716.4]
  wire  _T_6780; // @[OneHot.scala 66:30:@3717.4]
  wire  _T_6781; // @[OneHot.scala 66:30:@3718.4]
  wire  _T_6782; // @[OneHot.scala 66:30:@3719.4]
  wire  _T_6783; // @[OneHot.scala 66:30:@3720.4]
  wire  _T_6784; // @[OneHot.scala 66:30:@3721.4]
  wire  _T_6785; // @[OneHot.scala 66:30:@3722.4]
  wire  _T_6786; // @[OneHot.scala 66:30:@3723.4]
  wire  _T_6787; // @[OneHot.scala 66:30:@3724.4]
  wire  _T_6788; // @[OneHot.scala 66:30:@3725.4]
  wire  _T_6789; // @[OneHot.scala 66:30:@3726.4]
  wire  _T_6790; // @[OneHot.scala 66:30:@3727.4]
  wire  _T_6791; // @[OneHot.scala 66:30:@3728.4]
  wire  _T_6792; // @[OneHot.scala 66:30:@3729.4]
  wire  _T_6793; // @[OneHot.scala 66:30:@3730.4]
  wire  _T_6794; // @[OneHot.scala 66:30:@3731.4]
  wire [15:0] _T_6835; // @[Mux.scala 31:69:@3749.4]
  wire [15:0] _T_6836; // @[Mux.scala 31:69:@3750.4]
  wire [15:0] _T_6837; // @[Mux.scala 31:69:@3751.4]
  wire [15:0] _T_6838; // @[Mux.scala 31:69:@3752.4]
  wire [15:0] _T_6839; // @[Mux.scala 31:69:@3753.4]
  wire [15:0] _T_6840; // @[Mux.scala 31:69:@3754.4]
  wire [15:0] _T_6841; // @[Mux.scala 31:69:@3755.4]
  wire [15:0] _T_6842; // @[Mux.scala 31:69:@3756.4]
  wire [15:0] _T_6843; // @[Mux.scala 31:69:@3757.4]
  wire [15:0] _T_6844; // @[Mux.scala 31:69:@3758.4]
  wire [15:0] _T_6845; // @[Mux.scala 31:69:@3759.4]
  wire [15:0] _T_6846; // @[Mux.scala 31:69:@3760.4]
  wire [15:0] _T_6847; // @[Mux.scala 31:69:@3761.4]
  wire [15:0] _T_6848; // @[Mux.scala 31:69:@3762.4]
  wire [15:0] _T_6849; // @[Mux.scala 31:69:@3763.4]
  wire [15:0] _T_6850; // @[Mux.scala 31:69:@3764.4]
  wire  _T_6851; // @[OneHot.scala 66:30:@3765.4]
  wire  _T_6852; // @[OneHot.scala 66:30:@3766.4]
  wire  _T_6853; // @[OneHot.scala 66:30:@3767.4]
  wire  _T_6854; // @[OneHot.scala 66:30:@3768.4]
  wire  _T_6855; // @[OneHot.scala 66:30:@3769.4]
  wire  _T_6856; // @[OneHot.scala 66:30:@3770.4]
  wire  _T_6857; // @[OneHot.scala 66:30:@3771.4]
  wire  _T_6858; // @[OneHot.scala 66:30:@3772.4]
  wire  _T_6859; // @[OneHot.scala 66:30:@3773.4]
  wire  _T_6860; // @[OneHot.scala 66:30:@3774.4]
  wire  _T_6861; // @[OneHot.scala 66:30:@3775.4]
  wire  _T_6862; // @[OneHot.scala 66:30:@3776.4]
  wire  _T_6863; // @[OneHot.scala 66:30:@3777.4]
  wire  _T_6864; // @[OneHot.scala 66:30:@3778.4]
  wire  _T_6865; // @[OneHot.scala 66:30:@3779.4]
  wire  _T_6866; // @[OneHot.scala 66:30:@3780.4]
  wire [15:0] _T_6907; // @[Mux.scala 31:69:@3798.4]
  wire [15:0] _T_6908; // @[Mux.scala 31:69:@3799.4]
  wire [15:0] _T_6909; // @[Mux.scala 31:69:@3800.4]
  wire [15:0] _T_6910; // @[Mux.scala 31:69:@3801.4]
  wire [15:0] _T_6911; // @[Mux.scala 31:69:@3802.4]
  wire [15:0] _T_6912; // @[Mux.scala 31:69:@3803.4]
  wire [15:0] _T_6913; // @[Mux.scala 31:69:@3804.4]
  wire [15:0] _T_6914; // @[Mux.scala 31:69:@3805.4]
  wire [15:0] _T_6915; // @[Mux.scala 31:69:@3806.4]
  wire [15:0] _T_6916; // @[Mux.scala 31:69:@3807.4]
  wire [15:0] _T_6917; // @[Mux.scala 31:69:@3808.4]
  wire [15:0] _T_6918; // @[Mux.scala 31:69:@3809.4]
  wire [15:0] _T_6919; // @[Mux.scala 31:69:@3810.4]
  wire [15:0] _T_6920; // @[Mux.scala 31:69:@3811.4]
  wire [15:0] _T_6921; // @[Mux.scala 31:69:@3812.4]
  wire [15:0] _T_6922; // @[Mux.scala 31:69:@3813.4]
  wire  _T_6923; // @[OneHot.scala 66:30:@3814.4]
  wire  _T_6924; // @[OneHot.scala 66:30:@3815.4]
  wire  _T_6925; // @[OneHot.scala 66:30:@3816.4]
  wire  _T_6926; // @[OneHot.scala 66:30:@3817.4]
  wire  _T_6927; // @[OneHot.scala 66:30:@3818.4]
  wire  _T_6928; // @[OneHot.scala 66:30:@3819.4]
  wire  _T_6929; // @[OneHot.scala 66:30:@3820.4]
  wire  _T_6930; // @[OneHot.scala 66:30:@3821.4]
  wire  _T_6931; // @[OneHot.scala 66:30:@3822.4]
  wire  _T_6932; // @[OneHot.scala 66:30:@3823.4]
  wire  _T_6933; // @[OneHot.scala 66:30:@3824.4]
  wire  _T_6934; // @[OneHot.scala 66:30:@3825.4]
  wire  _T_6935; // @[OneHot.scala 66:30:@3826.4]
  wire  _T_6936; // @[OneHot.scala 66:30:@3827.4]
  wire  _T_6937; // @[OneHot.scala 66:30:@3828.4]
  wire  _T_6938; // @[OneHot.scala 66:30:@3829.4]
  wire [15:0] _T_6979; // @[Mux.scala 31:69:@3847.4]
  wire [15:0] _T_6980; // @[Mux.scala 31:69:@3848.4]
  wire [15:0] _T_6981; // @[Mux.scala 31:69:@3849.4]
  wire [15:0] _T_6982; // @[Mux.scala 31:69:@3850.4]
  wire [15:0] _T_6983; // @[Mux.scala 31:69:@3851.4]
  wire [15:0] _T_6984; // @[Mux.scala 31:69:@3852.4]
  wire [15:0] _T_6985; // @[Mux.scala 31:69:@3853.4]
  wire [15:0] _T_6986; // @[Mux.scala 31:69:@3854.4]
  wire [15:0] _T_6987; // @[Mux.scala 31:69:@3855.4]
  wire [15:0] _T_6988; // @[Mux.scala 31:69:@3856.4]
  wire [15:0] _T_6989; // @[Mux.scala 31:69:@3857.4]
  wire [15:0] _T_6990; // @[Mux.scala 31:69:@3858.4]
  wire [15:0] _T_6991; // @[Mux.scala 31:69:@3859.4]
  wire [15:0] _T_6992; // @[Mux.scala 31:69:@3860.4]
  wire [15:0] _T_6993; // @[Mux.scala 31:69:@3861.4]
  wire [15:0] _T_6994; // @[Mux.scala 31:69:@3862.4]
  wire  _T_6995; // @[OneHot.scala 66:30:@3863.4]
  wire  _T_6996; // @[OneHot.scala 66:30:@3864.4]
  wire  _T_6997; // @[OneHot.scala 66:30:@3865.4]
  wire  _T_6998; // @[OneHot.scala 66:30:@3866.4]
  wire  _T_6999; // @[OneHot.scala 66:30:@3867.4]
  wire  _T_7000; // @[OneHot.scala 66:30:@3868.4]
  wire  _T_7001; // @[OneHot.scala 66:30:@3869.4]
  wire  _T_7002; // @[OneHot.scala 66:30:@3870.4]
  wire  _T_7003; // @[OneHot.scala 66:30:@3871.4]
  wire  _T_7004; // @[OneHot.scala 66:30:@3872.4]
  wire  _T_7005; // @[OneHot.scala 66:30:@3873.4]
  wire  _T_7006; // @[OneHot.scala 66:30:@3874.4]
  wire  _T_7007; // @[OneHot.scala 66:30:@3875.4]
  wire  _T_7008; // @[OneHot.scala 66:30:@3876.4]
  wire  _T_7009; // @[OneHot.scala 66:30:@3877.4]
  wire  _T_7010; // @[OneHot.scala 66:30:@3878.4]
  wire [15:0] _T_7051; // @[Mux.scala 31:69:@3896.4]
  wire [15:0] _T_7052; // @[Mux.scala 31:69:@3897.4]
  wire [15:0] _T_7053; // @[Mux.scala 31:69:@3898.4]
  wire [15:0] _T_7054; // @[Mux.scala 31:69:@3899.4]
  wire [15:0] _T_7055; // @[Mux.scala 31:69:@3900.4]
  wire [15:0] _T_7056; // @[Mux.scala 31:69:@3901.4]
  wire [15:0] _T_7057; // @[Mux.scala 31:69:@3902.4]
  wire [15:0] _T_7058; // @[Mux.scala 31:69:@3903.4]
  wire [15:0] _T_7059; // @[Mux.scala 31:69:@3904.4]
  wire [15:0] _T_7060; // @[Mux.scala 31:69:@3905.4]
  wire [15:0] _T_7061; // @[Mux.scala 31:69:@3906.4]
  wire [15:0] _T_7062; // @[Mux.scala 31:69:@3907.4]
  wire [15:0] _T_7063; // @[Mux.scala 31:69:@3908.4]
  wire [15:0] _T_7064; // @[Mux.scala 31:69:@3909.4]
  wire [15:0] _T_7065; // @[Mux.scala 31:69:@3910.4]
  wire [15:0] _T_7066; // @[Mux.scala 31:69:@3911.4]
  wire  _T_7067; // @[OneHot.scala 66:30:@3912.4]
  wire  _T_7068; // @[OneHot.scala 66:30:@3913.4]
  wire  _T_7069; // @[OneHot.scala 66:30:@3914.4]
  wire  _T_7070; // @[OneHot.scala 66:30:@3915.4]
  wire  _T_7071; // @[OneHot.scala 66:30:@3916.4]
  wire  _T_7072; // @[OneHot.scala 66:30:@3917.4]
  wire  _T_7073; // @[OneHot.scala 66:30:@3918.4]
  wire  _T_7074; // @[OneHot.scala 66:30:@3919.4]
  wire  _T_7075; // @[OneHot.scala 66:30:@3920.4]
  wire  _T_7076; // @[OneHot.scala 66:30:@3921.4]
  wire  _T_7077; // @[OneHot.scala 66:30:@3922.4]
  wire  _T_7078; // @[OneHot.scala 66:30:@3923.4]
  wire  _T_7079; // @[OneHot.scala 66:30:@3924.4]
  wire  _T_7080; // @[OneHot.scala 66:30:@3925.4]
  wire  _T_7081; // @[OneHot.scala 66:30:@3926.4]
  wire  _T_7082; // @[OneHot.scala 66:30:@3927.4]
  wire [7:0] _T_7147; // @[Mux.scala 19:72:@3951.4]
  wire [15:0] _T_7155; // @[Mux.scala 19:72:@3959.4]
  wire [15:0] _T_7157; // @[Mux.scala 19:72:@3960.4]
  wire [7:0] _T_7164; // @[Mux.scala 19:72:@3967.4]
  wire [15:0] _T_7172; // @[Mux.scala 19:72:@3975.4]
  wire [15:0] _T_7174; // @[Mux.scala 19:72:@3976.4]
  wire [7:0] _T_7181; // @[Mux.scala 19:72:@3983.4]
  wire [15:0] _T_7189; // @[Mux.scala 19:72:@3991.4]
  wire [15:0] _T_7191; // @[Mux.scala 19:72:@3992.4]
  wire [7:0] _T_7198; // @[Mux.scala 19:72:@3999.4]
  wire [15:0] _T_7206; // @[Mux.scala 19:72:@4007.4]
  wire [15:0] _T_7208; // @[Mux.scala 19:72:@4008.4]
  wire [7:0] _T_7215; // @[Mux.scala 19:72:@4015.4]
  wire [15:0] _T_7223; // @[Mux.scala 19:72:@4023.4]
  wire [15:0] _T_7225; // @[Mux.scala 19:72:@4024.4]
  wire [7:0] _T_7232; // @[Mux.scala 19:72:@4031.4]
  wire [15:0] _T_7240; // @[Mux.scala 19:72:@4039.4]
  wire [15:0] _T_7242; // @[Mux.scala 19:72:@4040.4]
  wire [7:0] _T_7249; // @[Mux.scala 19:72:@4047.4]
  wire [15:0] _T_7257; // @[Mux.scala 19:72:@4055.4]
  wire [15:0] _T_7259; // @[Mux.scala 19:72:@4056.4]
  wire [7:0] _T_7266; // @[Mux.scala 19:72:@4063.4]
  wire [15:0] _T_7274; // @[Mux.scala 19:72:@4071.4]
  wire [15:0] _T_7276; // @[Mux.scala 19:72:@4072.4]
  wire [7:0] _T_7283; // @[Mux.scala 19:72:@4079.4]
  wire [15:0] _T_7291; // @[Mux.scala 19:72:@4087.4]
  wire [15:0] _T_7293; // @[Mux.scala 19:72:@4088.4]
  wire [7:0] _T_7300; // @[Mux.scala 19:72:@4095.4]
  wire [15:0] _T_7308; // @[Mux.scala 19:72:@4103.4]
  wire [15:0] _T_7310; // @[Mux.scala 19:72:@4104.4]
  wire [7:0] _T_7317; // @[Mux.scala 19:72:@4111.4]
  wire [15:0] _T_7325; // @[Mux.scala 19:72:@4119.4]
  wire [15:0] _T_7327; // @[Mux.scala 19:72:@4120.4]
  wire [7:0] _T_7334; // @[Mux.scala 19:72:@4127.4]
  wire [15:0] _T_7342; // @[Mux.scala 19:72:@4135.4]
  wire [15:0] _T_7344; // @[Mux.scala 19:72:@4136.4]
  wire [7:0] _T_7351; // @[Mux.scala 19:72:@4143.4]
  wire [15:0] _T_7359; // @[Mux.scala 19:72:@4151.4]
  wire [15:0] _T_7361; // @[Mux.scala 19:72:@4152.4]
  wire [7:0] _T_7368; // @[Mux.scala 19:72:@4159.4]
  wire [15:0] _T_7376; // @[Mux.scala 19:72:@4167.4]
  wire [15:0] _T_7378; // @[Mux.scala 19:72:@4168.4]
  wire [7:0] _T_7385; // @[Mux.scala 19:72:@4175.4]
  wire [15:0] _T_7393; // @[Mux.scala 19:72:@4183.4]
  wire [15:0] _T_7395; // @[Mux.scala 19:72:@4184.4]
  wire [7:0] _T_7402; // @[Mux.scala 19:72:@4191.4]
  wire [15:0] _T_7410; // @[Mux.scala 19:72:@4199.4]
  wire [15:0] _T_7412; // @[Mux.scala 19:72:@4200.4]
  wire [15:0] _T_7413; // @[Mux.scala 19:72:@4201.4]
  wire [15:0] _T_7414; // @[Mux.scala 19:72:@4202.4]
  wire [15:0] _T_7415; // @[Mux.scala 19:72:@4203.4]
  wire [15:0] _T_7416; // @[Mux.scala 19:72:@4204.4]
  wire [15:0] _T_7417; // @[Mux.scala 19:72:@4205.4]
  wire [15:0] _T_7418; // @[Mux.scala 19:72:@4206.4]
  wire [15:0] _T_7419; // @[Mux.scala 19:72:@4207.4]
  wire [15:0] _T_7420; // @[Mux.scala 19:72:@4208.4]
  wire [15:0] _T_7421; // @[Mux.scala 19:72:@4209.4]
  wire [15:0] _T_7422; // @[Mux.scala 19:72:@4210.4]
  wire [15:0] _T_7423; // @[Mux.scala 19:72:@4211.4]
  wire [15:0] _T_7424; // @[Mux.scala 19:72:@4212.4]
  wire [15:0] _T_7425; // @[Mux.scala 19:72:@4213.4]
  wire [15:0] _T_7426; // @[Mux.scala 19:72:@4214.4]
  wire [15:0] _T_7427; // @[Mux.scala 19:72:@4215.4]
  wire  inputDataPriorityPorts_0_0; // @[Mux.scala 19:72:@4219.4]
  wire  inputDataPriorityPorts_0_1; // @[Mux.scala 19:72:@4221.4]
  wire  inputDataPriorityPorts_0_2; // @[Mux.scala 19:72:@4223.4]
  wire  inputDataPriorityPorts_0_3; // @[Mux.scala 19:72:@4225.4]
  wire  inputDataPriorityPorts_0_4; // @[Mux.scala 19:72:@4227.4]
  wire  inputDataPriorityPorts_0_5; // @[Mux.scala 19:72:@4229.4]
  wire  inputDataPriorityPorts_0_6; // @[Mux.scala 19:72:@4231.4]
  wire  inputDataPriorityPorts_0_7; // @[Mux.scala 19:72:@4233.4]
  wire  inputDataPriorityPorts_0_8; // @[Mux.scala 19:72:@4235.4]
  wire  inputDataPriorityPorts_0_9; // @[Mux.scala 19:72:@4237.4]
  wire  inputDataPriorityPorts_0_10; // @[Mux.scala 19:72:@4239.4]
  wire  inputDataPriorityPorts_0_11; // @[Mux.scala 19:72:@4241.4]
  wire  inputDataPriorityPorts_0_12; // @[Mux.scala 19:72:@4243.4]
  wire  inputDataPriorityPorts_0_13; // @[Mux.scala 19:72:@4245.4]
  wire  inputDataPriorityPorts_0_14; // @[Mux.scala 19:72:@4247.4]
  wire  inputDataPriorityPorts_0_15; // @[Mux.scala 19:72:@4249.4]
  wire  _T_7573; // @[AxiStoreQueue.scala 214:52:@4273.6]
  wire  _T_7574; // @[AxiStoreQueue.scala 214:81:@4274.6]
  wire [30:0] _GEN_992; // @[AxiStoreQueue.scala 215:40:@4278.6]
  wire  _GEN_993; // @[AxiStoreQueue.scala 215:40:@4278.6]
  wire  _T_7590; // @[AxiStoreQueue.scala 220:52:@4283.6]
  wire  _T_7591; // @[AxiStoreQueue.scala 220:81:@4284.6]
  wire [31:0] _GEN_994; // @[AxiStoreQueue.scala 221:40:@4288.6]
  wire  _GEN_995; // @[AxiStoreQueue.scala 221:40:@4288.6]
  wire  _GEN_996; // @[AxiStoreQueue.scala 209:35:@4267.4]
  wire  _GEN_997; // @[AxiStoreQueue.scala 209:35:@4267.4]
  wire [30:0] _GEN_998; // @[AxiStoreQueue.scala 209:35:@4267.4]
  wire [31:0] _GEN_999; // @[AxiStoreQueue.scala 209:35:@4267.4]
  wire  _T_7609; // @[AxiStoreQueue.scala 214:52:@4299.6]
  wire  _T_7610; // @[AxiStoreQueue.scala 214:81:@4300.6]
  wire [30:0] _GEN_1000; // @[AxiStoreQueue.scala 215:40:@4304.6]
  wire  _GEN_1001; // @[AxiStoreQueue.scala 215:40:@4304.6]
  wire  _T_7626; // @[AxiStoreQueue.scala 220:52:@4309.6]
  wire  _T_7627; // @[AxiStoreQueue.scala 220:81:@4310.6]
  wire [31:0] _GEN_1002; // @[AxiStoreQueue.scala 221:40:@4314.6]
  wire  _GEN_1003; // @[AxiStoreQueue.scala 221:40:@4314.6]
  wire  _GEN_1004; // @[AxiStoreQueue.scala 209:35:@4293.4]
  wire  _GEN_1005; // @[AxiStoreQueue.scala 209:35:@4293.4]
  wire [30:0] _GEN_1006; // @[AxiStoreQueue.scala 209:35:@4293.4]
  wire [31:0] _GEN_1007; // @[AxiStoreQueue.scala 209:35:@4293.4]
  wire  _T_7645; // @[AxiStoreQueue.scala 214:52:@4325.6]
  wire  _T_7646; // @[AxiStoreQueue.scala 214:81:@4326.6]
  wire [30:0] _GEN_1008; // @[AxiStoreQueue.scala 215:40:@4330.6]
  wire  _GEN_1009; // @[AxiStoreQueue.scala 215:40:@4330.6]
  wire  _T_7662; // @[AxiStoreQueue.scala 220:52:@4335.6]
  wire  _T_7663; // @[AxiStoreQueue.scala 220:81:@4336.6]
  wire [31:0] _GEN_1010; // @[AxiStoreQueue.scala 221:40:@4340.6]
  wire  _GEN_1011; // @[AxiStoreQueue.scala 221:40:@4340.6]
  wire  _GEN_1012; // @[AxiStoreQueue.scala 209:35:@4319.4]
  wire  _GEN_1013; // @[AxiStoreQueue.scala 209:35:@4319.4]
  wire [30:0] _GEN_1014; // @[AxiStoreQueue.scala 209:35:@4319.4]
  wire [31:0] _GEN_1015; // @[AxiStoreQueue.scala 209:35:@4319.4]
  wire  _T_7681; // @[AxiStoreQueue.scala 214:52:@4351.6]
  wire  _T_7682; // @[AxiStoreQueue.scala 214:81:@4352.6]
  wire [30:0] _GEN_1016; // @[AxiStoreQueue.scala 215:40:@4356.6]
  wire  _GEN_1017; // @[AxiStoreQueue.scala 215:40:@4356.6]
  wire  _T_7698; // @[AxiStoreQueue.scala 220:52:@4361.6]
  wire  _T_7699; // @[AxiStoreQueue.scala 220:81:@4362.6]
  wire [31:0] _GEN_1018; // @[AxiStoreQueue.scala 221:40:@4366.6]
  wire  _GEN_1019; // @[AxiStoreQueue.scala 221:40:@4366.6]
  wire  _GEN_1020; // @[AxiStoreQueue.scala 209:35:@4345.4]
  wire  _GEN_1021; // @[AxiStoreQueue.scala 209:35:@4345.4]
  wire [30:0] _GEN_1022; // @[AxiStoreQueue.scala 209:35:@4345.4]
  wire [31:0] _GEN_1023; // @[AxiStoreQueue.scala 209:35:@4345.4]
  wire  _T_7717; // @[AxiStoreQueue.scala 214:52:@4377.6]
  wire  _T_7718; // @[AxiStoreQueue.scala 214:81:@4378.6]
  wire [30:0] _GEN_1024; // @[AxiStoreQueue.scala 215:40:@4382.6]
  wire  _GEN_1025; // @[AxiStoreQueue.scala 215:40:@4382.6]
  wire  _T_7734; // @[AxiStoreQueue.scala 220:52:@4387.6]
  wire  _T_7735; // @[AxiStoreQueue.scala 220:81:@4388.6]
  wire [31:0] _GEN_1026; // @[AxiStoreQueue.scala 221:40:@4392.6]
  wire  _GEN_1027; // @[AxiStoreQueue.scala 221:40:@4392.6]
  wire  _GEN_1028; // @[AxiStoreQueue.scala 209:35:@4371.4]
  wire  _GEN_1029; // @[AxiStoreQueue.scala 209:35:@4371.4]
  wire [30:0] _GEN_1030; // @[AxiStoreQueue.scala 209:35:@4371.4]
  wire [31:0] _GEN_1031; // @[AxiStoreQueue.scala 209:35:@4371.4]
  wire  _T_7753; // @[AxiStoreQueue.scala 214:52:@4403.6]
  wire  _T_7754; // @[AxiStoreQueue.scala 214:81:@4404.6]
  wire [30:0] _GEN_1032; // @[AxiStoreQueue.scala 215:40:@4408.6]
  wire  _GEN_1033; // @[AxiStoreQueue.scala 215:40:@4408.6]
  wire  _T_7770; // @[AxiStoreQueue.scala 220:52:@4413.6]
  wire  _T_7771; // @[AxiStoreQueue.scala 220:81:@4414.6]
  wire [31:0] _GEN_1034; // @[AxiStoreQueue.scala 221:40:@4418.6]
  wire  _GEN_1035; // @[AxiStoreQueue.scala 221:40:@4418.6]
  wire  _GEN_1036; // @[AxiStoreQueue.scala 209:35:@4397.4]
  wire  _GEN_1037; // @[AxiStoreQueue.scala 209:35:@4397.4]
  wire [30:0] _GEN_1038; // @[AxiStoreQueue.scala 209:35:@4397.4]
  wire [31:0] _GEN_1039; // @[AxiStoreQueue.scala 209:35:@4397.4]
  wire  _T_7789; // @[AxiStoreQueue.scala 214:52:@4429.6]
  wire  _T_7790; // @[AxiStoreQueue.scala 214:81:@4430.6]
  wire [30:0] _GEN_1040; // @[AxiStoreQueue.scala 215:40:@4434.6]
  wire  _GEN_1041; // @[AxiStoreQueue.scala 215:40:@4434.6]
  wire  _T_7806; // @[AxiStoreQueue.scala 220:52:@4439.6]
  wire  _T_7807; // @[AxiStoreQueue.scala 220:81:@4440.6]
  wire [31:0] _GEN_1042; // @[AxiStoreQueue.scala 221:40:@4444.6]
  wire  _GEN_1043; // @[AxiStoreQueue.scala 221:40:@4444.6]
  wire  _GEN_1044; // @[AxiStoreQueue.scala 209:35:@4423.4]
  wire  _GEN_1045; // @[AxiStoreQueue.scala 209:35:@4423.4]
  wire [30:0] _GEN_1046; // @[AxiStoreQueue.scala 209:35:@4423.4]
  wire [31:0] _GEN_1047; // @[AxiStoreQueue.scala 209:35:@4423.4]
  wire  _T_7825; // @[AxiStoreQueue.scala 214:52:@4455.6]
  wire  _T_7826; // @[AxiStoreQueue.scala 214:81:@4456.6]
  wire [30:0] _GEN_1048; // @[AxiStoreQueue.scala 215:40:@4460.6]
  wire  _GEN_1049; // @[AxiStoreQueue.scala 215:40:@4460.6]
  wire  _T_7842; // @[AxiStoreQueue.scala 220:52:@4465.6]
  wire  _T_7843; // @[AxiStoreQueue.scala 220:81:@4466.6]
  wire [31:0] _GEN_1050; // @[AxiStoreQueue.scala 221:40:@4470.6]
  wire  _GEN_1051; // @[AxiStoreQueue.scala 221:40:@4470.6]
  wire  _GEN_1052; // @[AxiStoreQueue.scala 209:35:@4449.4]
  wire  _GEN_1053; // @[AxiStoreQueue.scala 209:35:@4449.4]
  wire [30:0] _GEN_1054; // @[AxiStoreQueue.scala 209:35:@4449.4]
  wire [31:0] _GEN_1055; // @[AxiStoreQueue.scala 209:35:@4449.4]
  wire  _T_7861; // @[AxiStoreQueue.scala 214:52:@4481.6]
  wire  _T_7862; // @[AxiStoreQueue.scala 214:81:@4482.6]
  wire [30:0] _GEN_1056; // @[AxiStoreQueue.scala 215:40:@4486.6]
  wire  _GEN_1057; // @[AxiStoreQueue.scala 215:40:@4486.6]
  wire  _T_7878; // @[AxiStoreQueue.scala 220:52:@4491.6]
  wire  _T_7879; // @[AxiStoreQueue.scala 220:81:@4492.6]
  wire [31:0] _GEN_1058; // @[AxiStoreQueue.scala 221:40:@4496.6]
  wire  _GEN_1059; // @[AxiStoreQueue.scala 221:40:@4496.6]
  wire  _GEN_1060; // @[AxiStoreQueue.scala 209:35:@4475.4]
  wire  _GEN_1061; // @[AxiStoreQueue.scala 209:35:@4475.4]
  wire [30:0] _GEN_1062; // @[AxiStoreQueue.scala 209:35:@4475.4]
  wire [31:0] _GEN_1063; // @[AxiStoreQueue.scala 209:35:@4475.4]
  wire  _T_7897; // @[AxiStoreQueue.scala 214:52:@4507.6]
  wire  _T_7898; // @[AxiStoreQueue.scala 214:81:@4508.6]
  wire [30:0] _GEN_1064; // @[AxiStoreQueue.scala 215:40:@4512.6]
  wire  _GEN_1065; // @[AxiStoreQueue.scala 215:40:@4512.6]
  wire  _T_7914; // @[AxiStoreQueue.scala 220:52:@4517.6]
  wire  _T_7915; // @[AxiStoreQueue.scala 220:81:@4518.6]
  wire [31:0] _GEN_1066; // @[AxiStoreQueue.scala 221:40:@4522.6]
  wire  _GEN_1067; // @[AxiStoreQueue.scala 221:40:@4522.6]
  wire  _GEN_1068; // @[AxiStoreQueue.scala 209:35:@4501.4]
  wire  _GEN_1069; // @[AxiStoreQueue.scala 209:35:@4501.4]
  wire [30:0] _GEN_1070; // @[AxiStoreQueue.scala 209:35:@4501.4]
  wire [31:0] _GEN_1071; // @[AxiStoreQueue.scala 209:35:@4501.4]
  wire  _T_7933; // @[AxiStoreQueue.scala 214:52:@4533.6]
  wire  _T_7934; // @[AxiStoreQueue.scala 214:81:@4534.6]
  wire [30:0] _GEN_1072; // @[AxiStoreQueue.scala 215:40:@4538.6]
  wire  _GEN_1073; // @[AxiStoreQueue.scala 215:40:@4538.6]
  wire  _T_7950; // @[AxiStoreQueue.scala 220:52:@4543.6]
  wire  _T_7951; // @[AxiStoreQueue.scala 220:81:@4544.6]
  wire [31:0] _GEN_1074; // @[AxiStoreQueue.scala 221:40:@4548.6]
  wire  _GEN_1075; // @[AxiStoreQueue.scala 221:40:@4548.6]
  wire  _GEN_1076; // @[AxiStoreQueue.scala 209:35:@4527.4]
  wire  _GEN_1077; // @[AxiStoreQueue.scala 209:35:@4527.4]
  wire [30:0] _GEN_1078; // @[AxiStoreQueue.scala 209:35:@4527.4]
  wire [31:0] _GEN_1079; // @[AxiStoreQueue.scala 209:35:@4527.4]
  wire  _T_7969; // @[AxiStoreQueue.scala 214:52:@4559.6]
  wire  _T_7970; // @[AxiStoreQueue.scala 214:81:@4560.6]
  wire [30:0] _GEN_1080; // @[AxiStoreQueue.scala 215:40:@4564.6]
  wire  _GEN_1081; // @[AxiStoreQueue.scala 215:40:@4564.6]
  wire  _T_7986; // @[AxiStoreQueue.scala 220:52:@4569.6]
  wire  _T_7987; // @[AxiStoreQueue.scala 220:81:@4570.6]
  wire [31:0] _GEN_1082; // @[AxiStoreQueue.scala 221:40:@4574.6]
  wire  _GEN_1083; // @[AxiStoreQueue.scala 221:40:@4574.6]
  wire  _GEN_1084; // @[AxiStoreQueue.scala 209:35:@4553.4]
  wire  _GEN_1085; // @[AxiStoreQueue.scala 209:35:@4553.4]
  wire [30:0] _GEN_1086; // @[AxiStoreQueue.scala 209:35:@4553.4]
  wire [31:0] _GEN_1087; // @[AxiStoreQueue.scala 209:35:@4553.4]
  wire  _T_8005; // @[AxiStoreQueue.scala 214:52:@4585.6]
  wire  _T_8006; // @[AxiStoreQueue.scala 214:81:@4586.6]
  wire [30:0] _GEN_1088; // @[AxiStoreQueue.scala 215:40:@4590.6]
  wire  _GEN_1089; // @[AxiStoreQueue.scala 215:40:@4590.6]
  wire  _T_8022; // @[AxiStoreQueue.scala 220:52:@4595.6]
  wire  _T_8023; // @[AxiStoreQueue.scala 220:81:@4596.6]
  wire [31:0] _GEN_1090; // @[AxiStoreQueue.scala 221:40:@4600.6]
  wire  _GEN_1091; // @[AxiStoreQueue.scala 221:40:@4600.6]
  wire  _GEN_1092; // @[AxiStoreQueue.scala 209:35:@4579.4]
  wire  _GEN_1093; // @[AxiStoreQueue.scala 209:35:@4579.4]
  wire [30:0] _GEN_1094; // @[AxiStoreQueue.scala 209:35:@4579.4]
  wire [31:0] _GEN_1095; // @[AxiStoreQueue.scala 209:35:@4579.4]
  wire  _T_8041; // @[AxiStoreQueue.scala 214:52:@4611.6]
  wire  _T_8042; // @[AxiStoreQueue.scala 214:81:@4612.6]
  wire [30:0] _GEN_1096; // @[AxiStoreQueue.scala 215:40:@4616.6]
  wire  _GEN_1097; // @[AxiStoreQueue.scala 215:40:@4616.6]
  wire  _T_8058; // @[AxiStoreQueue.scala 220:52:@4621.6]
  wire  _T_8059; // @[AxiStoreQueue.scala 220:81:@4622.6]
  wire [31:0] _GEN_1098; // @[AxiStoreQueue.scala 221:40:@4626.6]
  wire  _GEN_1099; // @[AxiStoreQueue.scala 221:40:@4626.6]
  wire  _GEN_1100; // @[AxiStoreQueue.scala 209:35:@4605.4]
  wire  _GEN_1101; // @[AxiStoreQueue.scala 209:35:@4605.4]
  wire [30:0] _GEN_1102; // @[AxiStoreQueue.scala 209:35:@4605.4]
  wire [31:0] _GEN_1103; // @[AxiStoreQueue.scala 209:35:@4605.4]
  wire  _T_8077; // @[AxiStoreQueue.scala 214:52:@4637.6]
  wire  _T_8078; // @[AxiStoreQueue.scala 214:81:@4638.6]
  wire [30:0] _GEN_1104; // @[AxiStoreQueue.scala 215:40:@4642.6]
  wire  _GEN_1105; // @[AxiStoreQueue.scala 215:40:@4642.6]
  wire  _T_8094; // @[AxiStoreQueue.scala 220:52:@4647.6]
  wire  _T_8095; // @[AxiStoreQueue.scala 220:81:@4648.6]
  wire [31:0] _GEN_1106; // @[AxiStoreQueue.scala 221:40:@4652.6]
  wire  _GEN_1107; // @[AxiStoreQueue.scala 221:40:@4652.6]
  wire  _GEN_1108; // @[AxiStoreQueue.scala 209:35:@4631.4]
  wire  _GEN_1109; // @[AxiStoreQueue.scala 209:35:@4631.4]
  wire [30:0] _GEN_1110; // @[AxiStoreQueue.scala 209:35:@4631.4]
  wire [31:0] _GEN_1111; // @[AxiStoreQueue.scala 209:35:@4631.4]
  wire  _T_8113; // @[AxiStoreQueue.scala 214:52:@4663.6]
  wire  _T_8114; // @[AxiStoreQueue.scala 214:81:@4664.6]
  wire [30:0] _GEN_1112; // @[AxiStoreQueue.scala 215:40:@4668.6]
  wire  _GEN_1113; // @[AxiStoreQueue.scala 215:40:@4668.6]
  wire  _T_8130; // @[AxiStoreQueue.scala 220:52:@4673.6]
  wire  _T_8131; // @[AxiStoreQueue.scala 220:81:@4674.6]
  wire [31:0] _GEN_1114; // @[AxiStoreQueue.scala 221:40:@4678.6]
  wire  _GEN_1115; // @[AxiStoreQueue.scala 221:40:@4678.6]
  wire  _GEN_1116; // @[AxiStoreQueue.scala 209:35:@4657.4]
  wire  _GEN_1117; // @[AxiStoreQueue.scala 209:35:@4657.4]
  wire [30:0] _GEN_1118; // @[AxiStoreQueue.scala 209:35:@4657.4]
  wire [31:0] _GEN_1119; // @[AxiStoreQueue.scala 209:35:@4657.4]
  wire  _T_8145; // @[AxiStoreQueue.scala 234:30:@4683.4]
  wire [4:0] _T_8148; // @[util.scala 10:8:@4685.6]
  wire [4:0] _GEN_64; // @[util.scala 10:14:@4686.6]
  wire [4:0] _T_8149; // @[util.scala 10:14:@4686.6]
  wire [4:0] _GEN_1120; // @[AxiStoreQueue.scala 234:47:@4684.4]
  wire [3:0] _GEN_1251; // @[util.scala 10:8:@4698.6]
  wire [4:0] _T_8161; // @[util.scala 10:8:@4698.6]
  wire [4:0] _GEN_65; // @[util.scala 10:14:@4699.6]
  wire [4:0] _T_8162; // @[util.scala 10:14:@4699.6]
  wire [4:0] _GEN_1138; // @[AxiStoreQueue.scala 243:20:@4697.4]
  wire  _T_8164; // @[AxiStoreQueue.scala 247:84:@4702.4]
  wire  _T_8165; // @[AxiStoreQueue.scala 247:81:@4703.4]
  wire  _T_8167; // @[AxiStoreQueue.scala 247:84:@4704.4]
  wire  _T_8168; // @[AxiStoreQueue.scala 247:81:@4705.4]
  wire  _T_8170; // @[AxiStoreQueue.scala 247:84:@4706.4]
  wire  _T_8171; // @[AxiStoreQueue.scala 247:81:@4707.4]
  wire  _T_8173; // @[AxiStoreQueue.scala 247:84:@4708.4]
  wire  _T_8174; // @[AxiStoreQueue.scala 247:81:@4709.4]
  wire  _T_8176; // @[AxiStoreQueue.scala 247:84:@4710.4]
  wire  _T_8177; // @[AxiStoreQueue.scala 247:81:@4711.4]
  wire  _T_8179; // @[AxiStoreQueue.scala 247:84:@4712.4]
  wire  _T_8180; // @[AxiStoreQueue.scala 247:81:@4713.4]
  wire  _T_8182; // @[AxiStoreQueue.scala 247:84:@4714.4]
  wire  _T_8183; // @[AxiStoreQueue.scala 247:81:@4715.4]
  wire  _T_8185; // @[AxiStoreQueue.scala 247:84:@4716.4]
  wire  _T_8186; // @[AxiStoreQueue.scala 247:81:@4717.4]
  wire  _T_8188; // @[AxiStoreQueue.scala 247:84:@4718.4]
  wire  _T_8189; // @[AxiStoreQueue.scala 247:81:@4719.4]
  wire  _T_8191; // @[AxiStoreQueue.scala 247:84:@4720.4]
  wire  _T_8192; // @[AxiStoreQueue.scala 247:81:@4721.4]
  wire  _T_8194; // @[AxiStoreQueue.scala 247:84:@4722.4]
  wire  _T_8195; // @[AxiStoreQueue.scala 247:81:@4723.4]
  wire  _T_8197; // @[AxiStoreQueue.scala 247:84:@4724.4]
  wire  _T_8198; // @[AxiStoreQueue.scala 247:81:@4725.4]
  wire  _T_8200; // @[AxiStoreQueue.scala 247:84:@4726.4]
  wire  _T_8201; // @[AxiStoreQueue.scala 247:81:@4727.4]
  wire  _T_8203; // @[AxiStoreQueue.scala 247:84:@4728.4]
  wire  _T_8204; // @[AxiStoreQueue.scala 247:81:@4729.4]
  wire  _T_8206; // @[AxiStoreQueue.scala 247:84:@4730.4]
  wire  _T_8207; // @[AxiStoreQueue.scala 247:81:@4731.4]
  wire  _T_8209; // @[AxiStoreQueue.scala 247:84:@4732.4]
  wire  _T_8210; // @[AxiStoreQueue.scala 247:81:@4733.4]
  wire  _T_8235; // @[AxiStoreQueue.scala 247:98:@4752.4]
  wire  _T_8236; // @[AxiStoreQueue.scala 247:98:@4753.4]
  wire  _T_8237; // @[AxiStoreQueue.scala 247:98:@4754.4]
  wire  _T_8238; // @[AxiStoreQueue.scala 247:98:@4755.4]
  wire  _T_8239; // @[AxiStoreQueue.scala 247:98:@4756.4]
  wire  _T_8240; // @[AxiStoreQueue.scala 247:98:@4757.4]
  wire  _T_8241; // @[AxiStoreQueue.scala 247:98:@4758.4]
  wire  _T_8242; // @[AxiStoreQueue.scala 247:98:@4759.4]
  wire  _T_8243; // @[AxiStoreQueue.scala 247:98:@4760.4]
  wire  _T_8244; // @[AxiStoreQueue.scala 247:98:@4761.4]
  wire  _T_8245; // @[AxiStoreQueue.scala 247:98:@4762.4]
  wire  _T_8246; // @[AxiStoreQueue.scala 247:98:@4763.4]
  wire  _T_8247; // @[AxiStoreQueue.scala 247:98:@4764.4]
  wire  _T_8248; // @[AxiStoreQueue.scala 247:98:@4765.4]
  wire [31:0] _GEN_1140; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1141; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1142; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1143; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1144; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1145; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1146; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1147; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1148; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1149; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1150; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1151; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1152; // @[AxiStoreQueue.scala 262:21:@4835.4]
  wire [31:0] _GEN_1153; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1155 = {{2'd0}, tail}; // @[util.scala 14:20:@174.4]
  assign _T_1604 = 6'h10 - _GEN_1155; // @[util.scala 14:20:@174.4]
  assign _T_1605 = $unsigned(_T_1604); // @[util.scala 14:20:@175.4]
  assign _T_1606 = _T_1605[5:0]; // @[util.scala 14:20:@176.4]
  assign _GEN_0 = _T_1606 % 6'h10; // @[util.scala 14:25:@177.4]
  assign _T_1607 = _GEN_0[4:0]; // @[util.scala 14:25:@177.4]
  assign _GEN_1156 = {{4'd0}, io_bbNumStores}; // @[AxiStoreQueue.scala 72:46:@178.4]
  assign _T_1608 = _T_1607 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@178.4]
  assign initBits_0 = _T_1608 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@179.4]
  assign _T_1613 = 6'h11 - _GEN_1155; // @[util.scala 14:20:@181.4]
  assign _T_1614 = $unsigned(_T_1613); // @[util.scala 14:20:@182.4]
  assign _T_1615 = _T_1614[5:0]; // @[util.scala 14:20:@183.4]
  assign _GEN_16 = _T_1615 % 6'h10; // @[util.scala 14:25:@184.4]
  assign _T_1616 = _GEN_16[4:0]; // @[util.scala 14:25:@184.4]
  assign _T_1617 = _T_1616 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@185.4]
  assign initBits_1 = _T_1617 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@186.4]
  assign _T_1622 = 6'h12 - _GEN_1155; // @[util.scala 14:20:@188.4]
  assign _T_1623 = $unsigned(_T_1622); // @[util.scala 14:20:@189.4]
  assign _T_1624 = _T_1623[5:0]; // @[util.scala 14:20:@190.4]
  assign _GEN_17 = _T_1624 % 6'h10; // @[util.scala 14:25:@191.4]
  assign _T_1625 = _GEN_17[4:0]; // @[util.scala 14:25:@191.4]
  assign _T_1626 = _T_1625 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@192.4]
  assign initBits_2 = _T_1626 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@193.4]
  assign _T_1631 = 6'h13 - _GEN_1155; // @[util.scala 14:20:@195.4]
  assign _T_1632 = $unsigned(_T_1631); // @[util.scala 14:20:@196.4]
  assign _T_1633 = _T_1632[5:0]; // @[util.scala 14:20:@197.4]
  assign _GEN_18 = _T_1633 % 6'h10; // @[util.scala 14:25:@198.4]
  assign _T_1634 = _GEN_18[4:0]; // @[util.scala 14:25:@198.4]
  assign _T_1635 = _T_1634 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@199.4]
  assign initBits_3 = _T_1635 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@200.4]
  assign _T_1640 = 6'h14 - _GEN_1155; // @[util.scala 14:20:@202.4]
  assign _T_1641 = $unsigned(_T_1640); // @[util.scala 14:20:@203.4]
  assign _T_1642 = _T_1641[5:0]; // @[util.scala 14:20:@204.4]
  assign _GEN_19 = _T_1642 % 6'h10; // @[util.scala 14:25:@205.4]
  assign _T_1643 = _GEN_19[4:0]; // @[util.scala 14:25:@205.4]
  assign _T_1644 = _T_1643 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@206.4]
  assign initBits_4 = _T_1644 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@207.4]
  assign _T_1649 = 6'h15 - _GEN_1155; // @[util.scala 14:20:@209.4]
  assign _T_1650 = $unsigned(_T_1649); // @[util.scala 14:20:@210.4]
  assign _T_1651 = _T_1650[5:0]; // @[util.scala 14:20:@211.4]
  assign _GEN_20 = _T_1651 % 6'h10; // @[util.scala 14:25:@212.4]
  assign _T_1652 = _GEN_20[4:0]; // @[util.scala 14:25:@212.4]
  assign _T_1653 = _T_1652 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@213.4]
  assign initBits_5 = _T_1653 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@214.4]
  assign _T_1658 = 6'h16 - _GEN_1155; // @[util.scala 14:20:@216.4]
  assign _T_1659 = $unsigned(_T_1658); // @[util.scala 14:20:@217.4]
  assign _T_1660 = _T_1659[5:0]; // @[util.scala 14:20:@218.4]
  assign _GEN_21 = _T_1660 % 6'h10; // @[util.scala 14:25:@219.4]
  assign _T_1661 = _GEN_21[4:0]; // @[util.scala 14:25:@219.4]
  assign _T_1662 = _T_1661 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@220.4]
  assign initBits_6 = _T_1662 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@221.4]
  assign _T_1667 = 6'h17 - _GEN_1155; // @[util.scala 14:20:@223.4]
  assign _T_1668 = $unsigned(_T_1667); // @[util.scala 14:20:@224.4]
  assign _T_1669 = _T_1668[5:0]; // @[util.scala 14:20:@225.4]
  assign _GEN_22 = _T_1669 % 6'h10; // @[util.scala 14:25:@226.4]
  assign _T_1670 = _GEN_22[4:0]; // @[util.scala 14:25:@226.4]
  assign _T_1671 = _T_1670 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@227.4]
  assign initBits_7 = _T_1671 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@228.4]
  assign _T_1676 = 6'h18 - _GEN_1155; // @[util.scala 14:20:@230.4]
  assign _T_1677 = $unsigned(_T_1676); // @[util.scala 14:20:@231.4]
  assign _T_1678 = _T_1677[5:0]; // @[util.scala 14:20:@232.4]
  assign _GEN_23 = _T_1678 % 6'h10; // @[util.scala 14:25:@233.4]
  assign _T_1679 = _GEN_23[4:0]; // @[util.scala 14:25:@233.4]
  assign _T_1680 = _T_1679 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@234.4]
  assign initBits_8 = _T_1680 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@235.4]
  assign _T_1685 = 6'h19 - _GEN_1155; // @[util.scala 14:20:@237.4]
  assign _T_1686 = $unsigned(_T_1685); // @[util.scala 14:20:@238.4]
  assign _T_1687 = _T_1686[5:0]; // @[util.scala 14:20:@239.4]
  assign _GEN_24 = _T_1687 % 6'h10; // @[util.scala 14:25:@240.4]
  assign _T_1688 = _GEN_24[4:0]; // @[util.scala 14:25:@240.4]
  assign _T_1689 = _T_1688 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@241.4]
  assign initBits_9 = _T_1689 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@242.4]
  assign _T_1694 = 6'h1a - _GEN_1155; // @[util.scala 14:20:@244.4]
  assign _T_1695 = $unsigned(_T_1694); // @[util.scala 14:20:@245.4]
  assign _T_1696 = _T_1695[5:0]; // @[util.scala 14:20:@246.4]
  assign _GEN_25 = _T_1696 % 6'h10; // @[util.scala 14:25:@247.4]
  assign _T_1697 = _GEN_25[4:0]; // @[util.scala 14:25:@247.4]
  assign _T_1698 = _T_1697 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@248.4]
  assign initBits_10 = _T_1698 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@249.4]
  assign _T_1703 = 6'h1b - _GEN_1155; // @[util.scala 14:20:@251.4]
  assign _T_1704 = $unsigned(_T_1703); // @[util.scala 14:20:@252.4]
  assign _T_1705 = _T_1704[5:0]; // @[util.scala 14:20:@253.4]
  assign _GEN_26 = _T_1705 % 6'h10; // @[util.scala 14:25:@254.4]
  assign _T_1706 = _GEN_26[4:0]; // @[util.scala 14:25:@254.4]
  assign _T_1707 = _T_1706 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@255.4]
  assign initBits_11 = _T_1707 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@256.4]
  assign _T_1712 = 6'h1c - _GEN_1155; // @[util.scala 14:20:@258.4]
  assign _T_1713 = $unsigned(_T_1712); // @[util.scala 14:20:@259.4]
  assign _T_1714 = _T_1713[5:0]; // @[util.scala 14:20:@260.4]
  assign _GEN_27 = _T_1714 % 6'h10; // @[util.scala 14:25:@261.4]
  assign _T_1715 = _GEN_27[4:0]; // @[util.scala 14:25:@261.4]
  assign _T_1716 = _T_1715 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@262.4]
  assign initBits_12 = _T_1716 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@263.4]
  assign _T_1721 = 6'h1d - _GEN_1155; // @[util.scala 14:20:@265.4]
  assign _T_1722 = $unsigned(_T_1721); // @[util.scala 14:20:@266.4]
  assign _T_1723 = _T_1722[5:0]; // @[util.scala 14:20:@267.4]
  assign _GEN_28 = _T_1723 % 6'h10; // @[util.scala 14:25:@268.4]
  assign _T_1724 = _GEN_28[4:0]; // @[util.scala 14:25:@268.4]
  assign _T_1725 = _T_1724 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@269.4]
  assign initBits_13 = _T_1725 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@270.4]
  assign _T_1730 = 6'h1e - _GEN_1155; // @[util.scala 14:20:@272.4]
  assign _T_1731 = $unsigned(_T_1730); // @[util.scala 14:20:@273.4]
  assign _T_1732 = _T_1731[5:0]; // @[util.scala 14:20:@274.4]
  assign _GEN_29 = _T_1732 % 6'h10; // @[util.scala 14:25:@275.4]
  assign _T_1733 = _GEN_29[4:0]; // @[util.scala 14:25:@275.4]
  assign _T_1734 = _T_1733 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@276.4]
  assign initBits_14 = _T_1734 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@277.4]
  assign _T_1739 = 6'h1f - _GEN_1155; // @[util.scala 14:20:@279.4]
  assign _T_1740 = $unsigned(_T_1739); // @[util.scala 14:20:@280.4]
  assign _T_1741 = _T_1740[5:0]; // @[util.scala 14:20:@281.4]
  assign _GEN_30 = _T_1741 % 6'h10; // @[util.scala 14:25:@282.4]
  assign _T_1742 = _GEN_30[4:0]; // @[util.scala 14:25:@282.4]
  assign _T_1743 = _T_1742 < _GEN_1156; // @[AxiStoreQueue.scala 72:46:@283.4]
  assign initBits_15 = _T_1743 & io_bbStart; // @[AxiStoreQueue.scala 72:64:@284.4]
  assign _T_1766 = allocatedEntries_0 | initBits_0; // @[AxiStoreQueue.scala 74:78:@302.4]
  assign _T_1767 = allocatedEntries_1 | initBits_1; // @[AxiStoreQueue.scala 74:78:@303.4]
  assign _T_1768 = allocatedEntries_2 | initBits_2; // @[AxiStoreQueue.scala 74:78:@304.4]
  assign _T_1769 = allocatedEntries_3 | initBits_3; // @[AxiStoreQueue.scala 74:78:@305.4]
  assign _T_1770 = allocatedEntries_4 | initBits_4; // @[AxiStoreQueue.scala 74:78:@306.4]
  assign _T_1771 = allocatedEntries_5 | initBits_5; // @[AxiStoreQueue.scala 74:78:@307.4]
  assign _T_1772 = allocatedEntries_6 | initBits_6; // @[AxiStoreQueue.scala 74:78:@308.4]
  assign _T_1773 = allocatedEntries_7 | initBits_7; // @[AxiStoreQueue.scala 74:78:@309.4]
  assign _T_1774 = allocatedEntries_8 | initBits_8; // @[AxiStoreQueue.scala 74:78:@310.4]
  assign _T_1775 = allocatedEntries_9 | initBits_9; // @[AxiStoreQueue.scala 74:78:@311.4]
  assign _T_1776 = allocatedEntries_10 | initBits_10; // @[AxiStoreQueue.scala 74:78:@312.4]
  assign _T_1777 = allocatedEntries_11 | initBits_11; // @[AxiStoreQueue.scala 74:78:@313.4]
  assign _T_1778 = allocatedEntries_12 | initBits_12; // @[AxiStoreQueue.scala 74:78:@314.4]
  assign _T_1779 = allocatedEntries_13 | initBits_13; // @[AxiStoreQueue.scala 74:78:@315.4]
  assign _T_1780 = allocatedEntries_14 | initBits_14; // @[AxiStoreQueue.scala 74:78:@316.4]
  assign _T_1781 = allocatedEntries_15 | initBits_15; // @[AxiStoreQueue.scala 74:78:@317.4]
  assign _T_1812 = _T_1607[3:0]; // @[:@357.6]
  assign _GEN_1 = 4'h1 == _T_1812 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_2 = 4'h2 == _T_1812 ? io_bbStoreOffsets_2 : _GEN_1; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_3 = 4'h3 == _T_1812 ? io_bbStoreOffsets_3 : _GEN_2; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_4 = 4'h4 == _T_1812 ? io_bbStoreOffsets_4 : _GEN_3; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_5 = 4'h5 == _T_1812 ? io_bbStoreOffsets_5 : _GEN_4; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_6 = 4'h6 == _T_1812 ? io_bbStoreOffsets_6 : _GEN_5; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_7 = 4'h7 == _T_1812 ? io_bbStoreOffsets_7 : _GEN_6; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_8 = 4'h8 == _T_1812 ? io_bbStoreOffsets_8 : _GEN_7; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_9 = 4'h9 == _T_1812 ? io_bbStoreOffsets_9 : _GEN_8; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_10 = 4'ha == _T_1812 ? io_bbStoreOffsets_10 : _GEN_9; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_11 = 4'hb == _T_1812 ? io_bbStoreOffsets_11 : _GEN_10; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_12 = 4'hc == _T_1812 ? io_bbStoreOffsets_12 : _GEN_11; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_13 = 4'hd == _T_1812 ? io_bbStoreOffsets_13 : _GEN_12; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_14 = 4'he == _T_1812 ? io_bbStoreOffsets_14 : _GEN_13; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_15 = 4'hf == _T_1812 ? io_bbStoreOffsets_15 : _GEN_14; // @[AxiStoreQueue.scala 78:20:@358.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[AxiStoreQueue.scala 77:25:@351.4]
  assign _GEN_33 = initBits_0 ? 1'h0 : portQ_0; // @[AxiStoreQueue.scala 77:25:@351.4]
  assign _T_1830 = _T_1616[3:0]; // @[:@373.6]
  assign _GEN_35 = 4'h1 == _T_1830 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_36 = 4'h2 == _T_1830 ? io_bbStoreOffsets_2 : _GEN_35; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_37 = 4'h3 == _T_1830 ? io_bbStoreOffsets_3 : _GEN_36; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_38 = 4'h4 == _T_1830 ? io_bbStoreOffsets_4 : _GEN_37; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_39 = 4'h5 == _T_1830 ? io_bbStoreOffsets_5 : _GEN_38; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_40 = 4'h6 == _T_1830 ? io_bbStoreOffsets_6 : _GEN_39; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_41 = 4'h7 == _T_1830 ? io_bbStoreOffsets_7 : _GEN_40; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_42 = 4'h8 == _T_1830 ? io_bbStoreOffsets_8 : _GEN_41; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_43 = 4'h9 == _T_1830 ? io_bbStoreOffsets_9 : _GEN_42; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_44 = 4'ha == _T_1830 ? io_bbStoreOffsets_10 : _GEN_43; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_45 = 4'hb == _T_1830 ? io_bbStoreOffsets_11 : _GEN_44; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_46 = 4'hc == _T_1830 ? io_bbStoreOffsets_12 : _GEN_45; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_47 = 4'hd == _T_1830 ? io_bbStoreOffsets_13 : _GEN_46; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_48 = 4'he == _T_1830 ? io_bbStoreOffsets_14 : _GEN_47; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_49 = 4'hf == _T_1830 ? io_bbStoreOffsets_15 : _GEN_48; // @[AxiStoreQueue.scala 78:20:@374.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[AxiStoreQueue.scala 77:25:@367.4]
  assign _GEN_67 = initBits_1 ? 1'h0 : portQ_1; // @[AxiStoreQueue.scala 77:25:@367.4]
  assign _T_1848 = _T_1625[3:0]; // @[:@389.6]
  assign _GEN_69 = 4'h1 == _T_1848 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_70 = 4'h2 == _T_1848 ? io_bbStoreOffsets_2 : _GEN_69; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_71 = 4'h3 == _T_1848 ? io_bbStoreOffsets_3 : _GEN_70; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_72 = 4'h4 == _T_1848 ? io_bbStoreOffsets_4 : _GEN_71; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_73 = 4'h5 == _T_1848 ? io_bbStoreOffsets_5 : _GEN_72; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_74 = 4'h6 == _T_1848 ? io_bbStoreOffsets_6 : _GEN_73; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_75 = 4'h7 == _T_1848 ? io_bbStoreOffsets_7 : _GEN_74; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_76 = 4'h8 == _T_1848 ? io_bbStoreOffsets_8 : _GEN_75; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_77 = 4'h9 == _T_1848 ? io_bbStoreOffsets_9 : _GEN_76; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_78 = 4'ha == _T_1848 ? io_bbStoreOffsets_10 : _GEN_77; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_79 = 4'hb == _T_1848 ? io_bbStoreOffsets_11 : _GEN_78; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_80 = 4'hc == _T_1848 ? io_bbStoreOffsets_12 : _GEN_79; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_81 = 4'hd == _T_1848 ? io_bbStoreOffsets_13 : _GEN_80; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_82 = 4'he == _T_1848 ? io_bbStoreOffsets_14 : _GEN_81; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_83 = 4'hf == _T_1848 ? io_bbStoreOffsets_15 : _GEN_82; // @[AxiStoreQueue.scala 78:20:@390.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[AxiStoreQueue.scala 77:25:@383.4]
  assign _GEN_101 = initBits_2 ? 1'h0 : portQ_2; // @[AxiStoreQueue.scala 77:25:@383.4]
  assign _T_1866 = _T_1634[3:0]; // @[:@405.6]
  assign _GEN_103 = 4'h1 == _T_1866 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_104 = 4'h2 == _T_1866 ? io_bbStoreOffsets_2 : _GEN_103; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_105 = 4'h3 == _T_1866 ? io_bbStoreOffsets_3 : _GEN_104; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_106 = 4'h4 == _T_1866 ? io_bbStoreOffsets_4 : _GEN_105; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_107 = 4'h5 == _T_1866 ? io_bbStoreOffsets_5 : _GEN_106; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_108 = 4'h6 == _T_1866 ? io_bbStoreOffsets_6 : _GEN_107; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_109 = 4'h7 == _T_1866 ? io_bbStoreOffsets_7 : _GEN_108; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_110 = 4'h8 == _T_1866 ? io_bbStoreOffsets_8 : _GEN_109; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_111 = 4'h9 == _T_1866 ? io_bbStoreOffsets_9 : _GEN_110; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_112 = 4'ha == _T_1866 ? io_bbStoreOffsets_10 : _GEN_111; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_113 = 4'hb == _T_1866 ? io_bbStoreOffsets_11 : _GEN_112; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_114 = 4'hc == _T_1866 ? io_bbStoreOffsets_12 : _GEN_113; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_115 = 4'hd == _T_1866 ? io_bbStoreOffsets_13 : _GEN_114; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_116 = 4'he == _T_1866 ? io_bbStoreOffsets_14 : _GEN_115; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_117 = 4'hf == _T_1866 ? io_bbStoreOffsets_15 : _GEN_116; // @[AxiStoreQueue.scala 78:20:@406.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[AxiStoreQueue.scala 77:25:@399.4]
  assign _GEN_135 = initBits_3 ? 1'h0 : portQ_3; // @[AxiStoreQueue.scala 77:25:@399.4]
  assign _T_1884 = _T_1643[3:0]; // @[:@421.6]
  assign _GEN_137 = 4'h1 == _T_1884 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_138 = 4'h2 == _T_1884 ? io_bbStoreOffsets_2 : _GEN_137; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_139 = 4'h3 == _T_1884 ? io_bbStoreOffsets_3 : _GEN_138; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_140 = 4'h4 == _T_1884 ? io_bbStoreOffsets_4 : _GEN_139; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_141 = 4'h5 == _T_1884 ? io_bbStoreOffsets_5 : _GEN_140; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_142 = 4'h6 == _T_1884 ? io_bbStoreOffsets_6 : _GEN_141; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_143 = 4'h7 == _T_1884 ? io_bbStoreOffsets_7 : _GEN_142; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_144 = 4'h8 == _T_1884 ? io_bbStoreOffsets_8 : _GEN_143; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_145 = 4'h9 == _T_1884 ? io_bbStoreOffsets_9 : _GEN_144; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_146 = 4'ha == _T_1884 ? io_bbStoreOffsets_10 : _GEN_145; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_147 = 4'hb == _T_1884 ? io_bbStoreOffsets_11 : _GEN_146; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_148 = 4'hc == _T_1884 ? io_bbStoreOffsets_12 : _GEN_147; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_149 = 4'hd == _T_1884 ? io_bbStoreOffsets_13 : _GEN_148; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_150 = 4'he == _T_1884 ? io_bbStoreOffsets_14 : _GEN_149; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_151 = 4'hf == _T_1884 ? io_bbStoreOffsets_15 : _GEN_150; // @[AxiStoreQueue.scala 78:20:@422.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[AxiStoreQueue.scala 77:25:@415.4]
  assign _GEN_169 = initBits_4 ? 1'h0 : portQ_4; // @[AxiStoreQueue.scala 77:25:@415.4]
  assign _T_1902 = _T_1652[3:0]; // @[:@437.6]
  assign _GEN_171 = 4'h1 == _T_1902 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_172 = 4'h2 == _T_1902 ? io_bbStoreOffsets_2 : _GEN_171; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_173 = 4'h3 == _T_1902 ? io_bbStoreOffsets_3 : _GEN_172; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_174 = 4'h4 == _T_1902 ? io_bbStoreOffsets_4 : _GEN_173; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_175 = 4'h5 == _T_1902 ? io_bbStoreOffsets_5 : _GEN_174; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_176 = 4'h6 == _T_1902 ? io_bbStoreOffsets_6 : _GEN_175; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_177 = 4'h7 == _T_1902 ? io_bbStoreOffsets_7 : _GEN_176; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_178 = 4'h8 == _T_1902 ? io_bbStoreOffsets_8 : _GEN_177; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_179 = 4'h9 == _T_1902 ? io_bbStoreOffsets_9 : _GEN_178; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_180 = 4'ha == _T_1902 ? io_bbStoreOffsets_10 : _GEN_179; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_181 = 4'hb == _T_1902 ? io_bbStoreOffsets_11 : _GEN_180; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_182 = 4'hc == _T_1902 ? io_bbStoreOffsets_12 : _GEN_181; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_183 = 4'hd == _T_1902 ? io_bbStoreOffsets_13 : _GEN_182; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_184 = 4'he == _T_1902 ? io_bbStoreOffsets_14 : _GEN_183; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_185 = 4'hf == _T_1902 ? io_bbStoreOffsets_15 : _GEN_184; // @[AxiStoreQueue.scala 78:20:@438.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[AxiStoreQueue.scala 77:25:@431.4]
  assign _GEN_203 = initBits_5 ? 1'h0 : portQ_5; // @[AxiStoreQueue.scala 77:25:@431.4]
  assign _T_1920 = _T_1661[3:0]; // @[:@453.6]
  assign _GEN_205 = 4'h1 == _T_1920 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_206 = 4'h2 == _T_1920 ? io_bbStoreOffsets_2 : _GEN_205; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_207 = 4'h3 == _T_1920 ? io_bbStoreOffsets_3 : _GEN_206; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_208 = 4'h4 == _T_1920 ? io_bbStoreOffsets_4 : _GEN_207; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_209 = 4'h5 == _T_1920 ? io_bbStoreOffsets_5 : _GEN_208; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_210 = 4'h6 == _T_1920 ? io_bbStoreOffsets_6 : _GEN_209; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_211 = 4'h7 == _T_1920 ? io_bbStoreOffsets_7 : _GEN_210; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_212 = 4'h8 == _T_1920 ? io_bbStoreOffsets_8 : _GEN_211; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_213 = 4'h9 == _T_1920 ? io_bbStoreOffsets_9 : _GEN_212; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_214 = 4'ha == _T_1920 ? io_bbStoreOffsets_10 : _GEN_213; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_215 = 4'hb == _T_1920 ? io_bbStoreOffsets_11 : _GEN_214; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_216 = 4'hc == _T_1920 ? io_bbStoreOffsets_12 : _GEN_215; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_217 = 4'hd == _T_1920 ? io_bbStoreOffsets_13 : _GEN_216; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_218 = 4'he == _T_1920 ? io_bbStoreOffsets_14 : _GEN_217; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_219 = 4'hf == _T_1920 ? io_bbStoreOffsets_15 : _GEN_218; // @[AxiStoreQueue.scala 78:20:@454.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[AxiStoreQueue.scala 77:25:@447.4]
  assign _GEN_237 = initBits_6 ? 1'h0 : portQ_6; // @[AxiStoreQueue.scala 77:25:@447.4]
  assign _T_1938 = _T_1670[3:0]; // @[:@469.6]
  assign _GEN_239 = 4'h1 == _T_1938 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_240 = 4'h2 == _T_1938 ? io_bbStoreOffsets_2 : _GEN_239; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_241 = 4'h3 == _T_1938 ? io_bbStoreOffsets_3 : _GEN_240; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_242 = 4'h4 == _T_1938 ? io_bbStoreOffsets_4 : _GEN_241; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_243 = 4'h5 == _T_1938 ? io_bbStoreOffsets_5 : _GEN_242; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_244 = 4'h6 == _T_1938 ? io_bbStoreOffsets_6 : _GEN_243; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_245 = 4'h7 == _T_1938 ? io_bbStoreOffsets_7 : _GEN_244; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_246 = 4'h8 == _T_1938 ? io_bbStoreOffsets_8 : _GEN_245; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_247 = 4'h9 == _T_1938 ? io_bbStoreOffsets_9 : _GEN_246; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_248 = 4'ha == _T_1938 ? io_bbStoreOffsets_10 : _GEN_247; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_249 = 4'hb == _T_1938 ? io_bbStoreOffsets_11 : _GEN_248; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_250 = 4'hc == _T_1938 ? io_bbStoreOffsets_12 : _GEN_249; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_251 = 4'hd == _T_1938 ? io_bbStoreOffsets_13 : _GEN_250; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_252 = 4'he == _T_1938 ? io_bbStoreOffsets_14 : _GEN_251; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_253 = 4'hf == _T_1938 ? io_bbStoreOffsets_15 : _GEN_252; // @[AxiStoreQueue.scala 78:20:@470.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[AxiStoreQueue.scala 77:25:@463.4]
  assign _GEN_271 = initBits_7 ? 1'h0 : portQ_7; // @[AxiStoreQueue.scala 77:25:@463.4]
  assign _T_1956 = _T_1679[3:0]; // @[:@485.6]
  assign _GEN_273 = 4'h1 == _T_1956 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_274 = 4'h2 == _T_1956 ? io_bbStoreOffsets_2 : _GEN_273; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_275 = 4'h3 == _T_1956 ? io_bbStoreOffsets_3 : _GEN_274; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_276 = 4'h4 == _T_1956 ? io_bbStoreOffsets_4 : _GEN_275; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_277 = 4'h5 == _T_1956 ? io_bbStoreOffsets_5 : _GEN_276; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_278 = 4'h6 == _T_1956 ? io_bbStoreOffsets_6 : _GEN_277; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_279 = 4'h7 == _T_1956 ? io_bbStoreOffsets_7 : _GEN_278; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_280 = 4'h8 == _T_1956 ? io_bbStoreOffsets_8 : _GEN_279; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_281 = 4'h9 == _T_1956 ? io_bbStoreOffsets_9 : _GEN_280; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_282 = 4'ha == _T_1956 ? io_bbStoreOffsets_10 : _GEN_281; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_283 = 4'hb == _T_1956 ? io_bbStoreOffsets_11 : _GEN_282; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_284 = 4'hc == _T_1956 ? io_bbStoreOffsets_12 : _GEN_283; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_285 = 4'hd == _T_1956 ? io_bbStoreOffsets_13 : _GEN_284; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_286 = 4'he == _T_1956 ? io_bbStoreOffsets_14 : _GEN_285; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_287 = 4'hf == _T_1956 ? io_bbStoreOffsets_15 : _GEN_286; // @[AxiStoreQueue.scala 78:20:@486.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[AxiStoreQueue.scala 77:25:@479.4]
  assign _GEN_305 = initBits_8 ? 1'h0 : portQ_8; // @[AxiStoreQueue.scala 77:25:@479.4]
  assign _T_1974 = _T_1688[3:0]; // @[:@501.6]
  assign _GEN_307 = 4'h1 == _T_1974 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_308 = 4'h2 == _T_1974 ? io_bbStoreOffsets_2 : _GEN_307; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_309 = 4'h3 == _T_1974 ? io_bbStoreOffsets_3 : _GEN_308; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_310 = 4'h4 == _T_1974 ? io_bbStoreOffsets_4 : _GEN_309; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_311 = 4'h5 == _T_1974 ? io_bbStoreOffsets_5 : _GEN_310; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_312 = 4'h6 == _T_1974 ? io_bbStoreOffsets_6 : _GEN_311; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_313 = 4'h7 == _T_1974 ? io_bbStoreOffsets_7 : _GEN_312; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_314 = 4'h8 == _T_1974 ? io_bbStoreOffsets_8 : _GEN_313; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_315 = 4'h9 == _T_1974 ? io_bbStoreOffsets_9 : _GEN_314; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_316 = 4'ha == _T_1974 ? io_bbStoreOffsets_10 : _GEN_315; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_317 = 4'hb == _T_1974 ? io_bbStoreOffsets_11 : _GEN_316; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_318 = 4'hc == _T_1974 ? io_bbStoreOffsets_12 : _GEN_317; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_319 = 4'hd == _T_1974 ? io_bbStoreOffsets_13 : _GEN_318; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_320 = 4'he == _T_1974 ? io_bbStoreOffsets_14 : _GEN_319; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_321 = 4'hf == _T_1974 ? io_bbStoreOffsets_15 : _GEN_320; // @[AxiStoreQueue.scala 78:20:@502.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[AxiStoreQueue.scala 77:25:@495.4]
  assign _GEN_339 = initBits_9 ? 1'h0 : portQ_9; // @[AxiStoreQueue.scala 77:25:@495.4]
  assign _T_1992 = _T_1697[3:0]; // @[:@517.6]
  assign _GEN_341 = 4'h1 == _T_1992 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_342 = 4'h2 == _T_1992 ? io_bbStoreOffsets_2 : _GEN_341; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_343 = 4'h3 == _T_1992 ? io_bbStoreOffsets_3 : _GEN_342; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_344 = 4'h4 == _T_1992 ? io_bbStoreOffsets_4 : _GEN_343; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_345 = 4'h5 == _T_1992 ? io_bbStoreOffsets_5 : _GEN_344; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_346 = 4'h6 == _T_1992 ? io_bbStoreOffsets_6 : _GEN_345; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_347 = 4'h7 == _T_1992 ? io_bbStoreOffsets_7 : _GEN_346; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_348 = 4'h8 == _T_1992 ? io_bbStoreOffsets_8 : _GEN_347; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_349 = 4'h9 == _T_1992 ? io_bbStoreOffsets_9 : _GEN_348; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_350 = 4'ha == _T_1992 ? io_bbStoreOffsets_10 : _GEN_349; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_351 = 4'hb == _T_1992 ? io_bbStoreOffsets_11 : _GEN_350; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_352 = 4'hc == _T_1992 ? io_bbStoreOffsets_12 : _GEN_351; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_353 = 4'hd == _T_1992 ? io_bbStoreOffsets_13 : _GEN_352; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_354 = 4'he == _T_1992 ? io_bbStoreOffsets_14 : _GEN_353; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_355 = 4'hf == _T_1992 ? io_bbStoreOffsets_15 : _GEN_354; // @[AxiStoreQueue.scala 78:20:@518.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[AxiStoreQueue.scala 77:25:@511.4]
  assign _GEN_373 = initBits_10 ? 1'h0 : portQ_10; // @[AxiStoreQueue.scala 77:25:@511.4]
  assign _T_2010 = _T_1706[3:0]; // @[:@533.6]
  assign _GEN_375 = 4'h1 == _T_2010 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_376 = 4'h2 == _T_2010 ? io_bbStoreOffsets_2 : _GEN_375; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_377 = 4'h3 == _T_2010 ? io_bbStoreOffsets_3 : _GEN_376; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_378 = 4'h4 == _T_2010 ? io_bbStoreOffsets_4 : _GEN_377; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_379 = 4'h5 == _T_2010 ? io_bbStoreOffsets_5 : _GEN_378; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_380 = 4'h6 == _T_2010 ? io_bbStoreOffsets_6 : _GEN_379; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_381 = 4'h7 == _T_2010 ? io_bbStoreOffsets_7 : _GEN_380; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_382 = 4'h8 == _T_2010 ? io_bbStoreOffsets_8 : _GEN_381; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_383 = 4'h9 == _T_2010 ? io_bbStoreOffsets_9 : _GEN_382; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_384 = 4'ha == _T_2010 ? io_bbStoreOffsets_10 : _GEN_383; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_385 = 4'hb == _T_2010 ? io_bbStoreOffsets_11 : _GEN_384; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_386 = 4'hc == _T_2010 ? io_bbStoreOffsets_12 : _GEN_385; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_387 = 4'hd == _T_2010 ? io_bbStoreOffsets_13 : _GEN_386; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_388 = 4'he == _T_2010 ? io_bbStoreOffsets_14 : _GEN_387; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_389 = 4'hf == _T_2010 ? io_bbStoreOffsets_15 : _GEN_388; // @[AxiStoreQueue.scala 78:20:@534.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[AxiStoreQueue.scala 77:25:@527.4]
  assign _GEN_407 = initBits_11 ? 1'h0 : portQ_11; // @[AxiStoreQueue.scala 77:25:@527.4]
  assign _T_2028 = _T_1715[3:0]; // @[:@549.6]
  assign _GEN_409 = 4'h1 == _T_2028 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_410 = 4'h2 == _T_2028 ? io_bbStoreOffsets_2 : _GEN_409; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_411 = 4'h3 == _T_2028 ? io_bbStoreOffsets_3 : _GEN_410; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_412 = 4'h4 == _T_2028 ? io_bbStoreOffsets_4 : _GEN_411; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_413 = 4'h5 == _T_2028 ? io_bbStoreOffsets_5 : _GEN_412; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_414 = 4'h6 == _T_2028 ? io_bbStoreOffsets_6 : _GEN_413; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_415 = 4'h7 == _T_2028 ? io_bbStoreOffsets_7 : _GEN_414; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_416 = 4'h8 == _T_2028 ? io_bbStoreOffsets_8 : _GEN_415; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_417 = 4'h9 == _T_2028 ? io_bbStoreOffsets_9 : _GEN_416; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_418 = 4'ha == _T_2028 ? io_bbStoreOffsets_10 : _GEN_417; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_419 = 4'hb == _T_2028 ? io_bbStoreOffsets_11 : _GEN_418; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_420 = 4'hc == _T_2028 ? io_bbStoreOffsets_12 : _GEN_419; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_421 = 4'hd == _T_2028 ? io_bbStoreOffsets_13 : _GEN_420; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_422 = 4'he == _T_2028 ? io_bbStoreOffsets_14 : _GEN_421; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_423 = 4'hf == _T_2028 ? io_bbStoreOffsets_15 : _GEN_422; // @[AxiStoreQueue.scala 78:20:@550.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[AxiStoreQueue.scala 77:25:@543.4]
  assign _GEN_441 = initBits_12 ? 1'h0 : portQ_12; // @[AxiStoreQueue.scala 77:25:@543.4]
  assign _T_2046 = _T_1724[3:0]; // @[:@565.6]
  assign _GEN_443 = 4'h1 == _T_2046 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_444 = 4'h2 == _T_2046 ? io_bbStoreOffsets_2 : _GEN_443; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_445 = 4'h3 == _T_2046 ? io_bbStoreOffsets_3 : _GEN_444; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_446 = 4'h4 == _T_2046 ? io_bbStoreOffsets_4 : _GEN_445; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_447 = 4'h5 == _T_2046 ? io_bbStoreOffsets_5 : _GEN_446; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_448 = 4'h6 == _T_2046 ? io_bbStoreOffsets_6 : _GEN_447; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_449 = 4'h7 == _T_2046 ? io_bbStoreOffsets_7 : _GEN_448; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_450 = 4'h8 == _T_2046 ? io_bbStoreOffsets_8 : _GEN_449; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_451 = 4'h9 == _T_2046 ? io_bbStoreOffsets_9 : _GEN_450; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_452 = 4'ha == _T_2046 ? io_bbStoreOffsets_10 : _GEN_451; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_453 = 4'hb == _T_2046 ? io_bbStoreOffsets_11 : _GEN_452; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_454 = 4'hc == _T_2046 ? io_bbStoreOffsets_12 : _GEN_453; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_455 = 4'hd == _T_2046 ? io_bbStoreOffsets_13 : _GEN_454; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_456 = 4'he == _T_2046 ? io_bbStoreOffsets_14 : _GEN_455; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_457 = 4'hf == _T_2046 ? io_bbStoreOffsets_15 : _GEN_456; // @[AxiStoreQueue.scala 78:20:@566.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[AxiStoreQueue.scala 77:25:@559.4]
  assign _GEN_475 = initBits_13 ? 1'h0 : portQ_13; // @[AxiStoreQueue.scala 77:25:@559.4]
  assign _T_2064 = _T_1733[3:0]; // @[:@581.6]
  assign _GEN_477 = 4'h1 == _T_2064 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_478 = 4'h2 == _T_2064 ? io_bbStoreOffsets_2 : _GEN_477; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_479 = 4'h3 == _T_2064 ? io_bbStoreOffsets_3 : _GEN_478; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_480 = 4'h4 == _T_2064 ? io_bbStoreOffsets_4 : _GEN_479; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_481 = 4'h5 == _T_2064 ? io_bbStoreOffsets_5 : _GEN_480; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_482 = 4'h6 == _T_2064 ? io_bbStoreOffsets_6 : _GEN_481; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_483 = 4'h7 == _T_2064 ? io_bbStoreOffsets_7 : _GEN_482; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_484 = 4'h8 == _T_2064 ? io_bbStoreOffsets_8 : _GEN_483; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_485 = 4'h9 == _T_2064 ? io_bbStoreOffsets_9 : _GEN_484; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_486 = 4'ha == _T_2064 ? io_bbStoreOffsets_10 : _GEN_485; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_487 = 4'hb == _T_2064 ? io_bbStoreOffsets_11 : _GEN_486; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_488 = 4'hc == _T_2064 ? io_bbStoreOffsets_12 : _GEN_487; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_489 = 4'hd == _T_2064 ? io_bbStoreOffsets_13 : _GEN_488; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_490 = 4'he == _T_2064 ? io_bbStoreOffsets_14 : _GEN_489; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_491 = 4'hf == _T_2064 ? io_bbStoreOffsets_15 : _GEN_490; // @[AxiStoreQueue.scala 78:20:@582.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[AxiStoreQueue.scala 77:25:@575.4]
  assign _GEN_509 = initBits_14 ? 1'h0 : portQ_14; // @[AxiStoreQueue.scala 77:25:@575.4]
  assign _T_2082 = _T_1742[3:0]; // @[:@597.6]
  assign _GEN_511 = 4'h1 == _T_2082 ? io_bbStoreOffsets_1 : io_bbStoreOffsets_0; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_512 = 4'h2 == _T_2082 ? io_bbStoreOffsets_2 : _GEN_511; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_513 = 4'h3 == _T_2082 ? io_bbStoreOffsets_3 : _GEN_512; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_514 = 4'h4 == _T_2082 ? io_bbStoreOffsets_4 : _GEN_513; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_515 = 4'h5 == _T_2082 ? io_bbStoreOffsets_5 : _GEN_514; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_516 = 4'h6 == _T_2082 ? io_bbStoreOffsets_6 : _GEN_515; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_517 = 4'h7 == _T_2082 ? io_bbStoreOffsets_7 : _GEN_516; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_518 = 4'h8 == _T_2082 ? io_bbStoreOffsets_8 : _GEN_517; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_519 = 4'h9 == _T_2082 ? io_bbStoreOffsets_9 : _GEN_518; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_520 = 4'ha == _T_2082 ? io_bbStoreOffsets_10 : _GEN_519; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_521 = 4'hb == _T_2082 ? io_bbStoreOffsets_11 : _GEN_520; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_522 = 4'hc == _T_2082 ? io_bbStoreOffsets_12 : _GEN_521; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_523 = 4'hd == _T_2082 ? io_bbStoreOffsets_13 : _GEN_522; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_524 = 4'he == _T_2082 ? io_bbStoreOffsets_14 : _GEN_523; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_525 = 4'hf == _T_2082 ? io_bbStoreOffsets_15 : _GEN_524; // @[AxiStoreQueue.scala 78:20:@598.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[AxiStoreQueue.scala 77:25:@591.4]
  assign _GEN_543 = initBits_15 ? 1'h0 : portQ_15; // @[AxiStoreQueue.scala 77:25:@591.4]
  assign _T_2104 = _GEN_15 + 4'h1; // @[util.scala 10:8:@616.6]
  assign _GEN_31 = _T_2104 % 5'h10; // @[util.scala 10:14:@617.6]
  assign _T_2105 = _GEN_31[4:0]; // @[util.scala 10:14:@617.6]
  assign _GEN_1220 = {{1'd0}, io_loadTail}; // @[AxiStoreQueue.scala 98:56:@618.6]
  assign _T_2106 = _T_2105 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@618.6]
  assign _T_2107 = io_loadEmpty & _T_2106; // @[AxiStoreQueue.scala 97:50:@619.6]
  assign _T_2109 = _T_2107 == 1'h0; // @[AxiStoreQueue.scala 97:35:@620.6]
  assign _T_2111 = previousLoadHead <= offsetQ_0; // @[AxiStoreQueue.scala 102:35:@628.8]
  assign _T_2112 = offsetQ_0 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@629.8]
  assign _T_2113 = _T_2111 & _T_2112; // @[AxiStoreQueue.scala 102:61:@630.8]
  assign _T_2115 = previousLoadHead > io_loadHead; // @[AxiStoreQueue.scala 104:35:@635.10]
  assign _T_2116 = io_loadHead <= offsetQ_0; // @[AxiStoreQueue.scala 105:23:@636.10]
  assign _T_2117 = offsetQ_0 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@637.10]
  assign _T_2118 = _T_2116 & _T_2117; // @[AxiStoreQueue.scala 105:49:@638.10]
  assign _T_2120 = _T_2118 == 1'h0; // @[AxiStoreQueue.scala 105:9:@639.10]
  assign _T_2121 = _T_2115 & _T_2120; // @[AxiStoreQueue.scala 104:49:@640.10]
  assign _GEN_560 = _T_2121 ? 1'h0 : checkBits_0; // @[AxiStoreQueue.scala 105:96:@641.10]
  assign _GEN_561 = _T_2113 ? 1'h0 : _GEN_560; // @[AxiStoreQueue.scala 102:102:@631.8]
  assign _GEN_562 = io_loadEmpty ? 1'h0 : _GEN_561; // @[AxiStoreQueue.scala 100:26:@624.6]
  assign _GEN_563 = initBits_0 ? _T_2109 : _GEN_562; // @[AxiStoreQueue.scala 96:35:@609.4]
  assign _T_2134 = _GEN_49 + 4'h1; // @[util.scala 10:8:@652.6]
  assign _GEN_34 = _T_2134 % 5'h10; // @[util.scala 10:14:@653.6]
  assign _T_2135 = _GEN_34[4:0]; // @[util.scala 10:14:@653.6]
  assign _T_2136 = _T_2135 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@654.6]
  assign _T_2137 = io_loadEmpty & _T_2136; // @[AxiStoreQueue.scala 97:50:@655.6]
  assign _T_2139 = _T_2137 == 1'h0; // @[AxiStoreQueue.scala 97:35:@656.6]
  assign _T_2141 = previousLoadHead <= offsetQ_1; // @[AxiStoreQueue.scala 102:35:@664.8]
  assign _T_2142 = offsetQ_1 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@665.8]
  assign _T_2143 = _T_2141 & _T_2142; // @[AxiStoreQueue.scala 102:61:@666.8]
  assign _T_2146 = io_loadHead <= offsetQ_1; // @[AxiStoreQueue.scala 105:23:@672.10]
  assign _T_2147 = offsetQ_1 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@673.10]
  assign _T_2148 = _T_2146 & _T_2147; // @[AxiStoreQueue.scala 105:49:@674.10]
  assign _T_2150 = _T_2148 == 1'h0; // @[AxiStoreQueue.scala 105:9:@675.10]
  assign _T_2151 = _T_2115 & _T_2150; // @[AxiStoreQueue.scala 104:49:@676.10]
  assign _GEN_580 = _T_2151 ? 1'h0 : checkBits_1; // @[AxiStoreQueue.scala 105:96:@677.10]
  assign _GEN_581 = _T_2143 ? 1'h0 : _GEN_580; // @[AxiStoreQueue.scala 102:102:@667.8]
  assign _GEN_582 = io_loadEmpty ? 1'h0 : _GEN_581; // @[AxiStoreQueue.scala 100:26:@660.6]
  assign _GEN_583 = initBits_1 ? _T_2139 : _GEN_582; // @[AxiStoreQueue.scala 96:35:@645.4]
  assign _T_2164 = _GEN_83 + 4'h1; // @[util.scala 10:8:@688.6]
  assign _GEN_50 = _T_2164 % 5'h10; // @[util.scala 10:14:@689.6]
  assign _T_2165 = _GEN_50[4:0]; // @[util.scala 10:14:@689.6]
  assign _T_2166 = _T_2165 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@690.6]
  assign _T_2167 = io_loadEmpty & _T_2166; // @[AxiStoreQueue.scala 97:50:@691.6]
  assign _T_2169 = _T_2167 == 1'h0; // @[AxiStoreQueue.scala 97:35:@692.6]
  assign _T_2171 = previousLoadHead <= offsetQ_2; // @[AxiStoreQueue.scala 102:35:@700.8]
  assign _T_2172 = offsetQ_2 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@701.8]
  assign _T_2173 = _T_2171 & _T_2172; // @[AxiStoreQueue.scala 102:61:@702.8]
  assign _T_2176 = io_loadHead <= offsetQ_2; // @[AxiStoreQueue.scala 105:23:@708.10]
  assign _T_2177 = offsetQ_2 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@709.10]
  assign _T_2178 = _T_2176 & _T_2177; // @[AxiStoreQueue.scala 105:49:@710.10]
  assign _T_2180 = _T_2178 == 1'h0; // @[AxiStoreQueue.scala 105:9:@711.10]
  assign _T_2181 = _T_2115 & _T_2180; // @[AxiStoreQueue.scala 104:49:@712.10]
  assign _GEN_600 = _T_2181 ? 1'h0 : checkBits_2; // @[AxiStoreQueue.scala 105:96:@713.10]
  assign _GEN_601 = _T_2173 ? 1'h0 : _GEN_600; // @[AxiStoreQueue.scala 102:102:@703.8]
  assign _GEN_602 = io_loadEmpty ? 1'h0 : _GEN_601; // @[AxiStoreQueue.scala 100:26:@696.6]
  assign _GEN_603 = initBits_2 ? _T_2169 : _GEN_602; // @[AxiStoreQueue.scala 96:35:@681.4]
  assign _T_2194 = _GEN_117 + 4'h1; // @[util.scala 10:8:@724.6]
  assign _GEN_51 = _T_2194 % 5'h10; // @[util.scala 10:14:@725.6]
  assign _T_2195 = _GEN_51[4:0]; // @[util.scala 10:14:@725.6]
  assign _T_2196 = _T_2195 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@726.6]
  assign _T_2197 = io_loadEmpty & _T_2196; // @[AxiStoreQueue.scala 97:50:@727.6]
  assign _T_2199 = _T_2197 == 1'h0; // @[AxiStoreQueue.scala 97:35:@728.6]
  assign _T_2201 = previousLoadHead <= offsetQ_3; // @[AxiStoreQueue.scala 102:35:@736.8]
  assign _T_2202 = offsetQ_3 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@737.8]
  assign _T_2203 = _T_2201 & _T_2202; // @[AxiStoreQueue.scala 102:61:@738.8]
  assign _T_2206 = io_loadHead <= offsetQ_3; // @[AxiStoreQueue.scala 105:23:@744.10]
  assign _T_2207 = offsetQ_3 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@745.10]
  assign _T_2208 = _T_2206 & _T_2207; // @[AxiStoreQueue.scala 105:49:@746.10]
  assign _T_2210 = _T_2208 == 1'h0; // @[AxiStoreQueue.scala 105:9:@747.10]
  assign _T_2211 = _T_2115 & _T_2210; // @[AxiStoreQueue.scala 104:49:@748.10]
  assign _GEN_620 = _T_2211 ? 1'h0 : checkBits_3; // @[AxiStoreQueue.scala 105:96:@749.10]
  assign _GEN_621 = _T_2203 ? 1'h0 : _GEN_620; // @[AxiStoreQueue.scala 102:102:@739.8]
  assign _GEN_622 = io_loadEmpty ? 1'h0 : _GEN_621; // @[AxiStoreQueue.scala 100:26:@732.6]
  assign _GEN_623 = initBits_3 ? _T_2199 : _GEN_622; // @[AxiStoreQueue.scala 96:35:@717.4]
  assign _T_2224 = _GEN_151 + 4'h1; // @[util.scala 10:8:@760.6]
  assign _GEN_52 = _T_2224 % 5'h10; // @[util.scala 10:14:@761.6]
  assign _T_2225 = _GEN_52[4:0]; // @[util.scala 10:14:@761.6]
  assign _T_2226 = _T_2225 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@762.6]
  assign _T_2227 = io_loadEmpty & _T_2226; // @[AxiStoreQueue.scala 97:50:@763.6]
  assign _T_2229 = _T_2227 == 1'h0; // @[AxiStoreQueue.scala 97:35:@764.6]
  assign _T_2231 = previousLoadHead <= offsetQ_4; // @[AxiStoreQueue.scala 102:35:@772.8]
  assign _T_2232 = offsetQ_4 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@773.8]
  assign _T_2233 = _T_2231 & _T_2232; // @[AxiStoreQueue.scala 102:61:@774.8]
  assign _T_2236 = io_loadHead <= offsetQ_4; // @[AxiStoreQueue.scala 105:23:@780.10]
  assign _T_2237 = offsetQ_4 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@781.10]
  assign _T_2238 = _T_2236 & _T_2237; // @[AxiStoreQueue.scala 105:49:@782.10]
  assign _T_2240 = _T_2238 == 1'h0; // @[AxiStoreQueue.scala 105:9:@783.10]
  assign _T_2241 = _T_2115 & _T_2240; // @[AxiStoreQueue.scala 104:49:@784.10]
  assign _GEN_640 = _T_2241 ? 1'h0 : checkBits_4; // @[AxiStoreQueue.scala 105:96:@785.10]
  assign _GEN_641 = _T_2233 ? 1'h0 : _GEN_640; // @[AxiStoreQueue.scala 102:102:@775.8]
  assign _GEN_642 = io_loadEmpty ? 1'h0 : _GEN_641; // @[AxiStoreQueue.scala 100:26:@768.6]
  assign _GEN_643 = initBits_4 ? _T_2229 : _GEN_642; // @[AxiStoreQueue.scala 96:35:@753.4]
  assign _T_2254 = _GEN_185 + 4'h1; // @[util.scala 10:8:@796.6]
  assign _GEN_53 = _T_2254 % 5'h10; // @[util.scala 10:14:@797.6]
  assign _T_2255 = _GEN_53[4:0]; // @[util.scala 10:14:@797.6]
  assign _T_2256 = _T_2255 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@798.6]
  assign _T_2257 = io_loadEmpty & _T_2256; // @[AxiStoreQueue.scala 97:50:@799.6]
  assign _T_2259 = _T_2257 == 1'h0; // @[AxiStoreQueue.scala 97:35:@800.6]
  assign _T_2261 = previousLoadHead <= offsetQ_5; // @[AxiStoreQueue.scala 102:35:@808.8]
  assign _T_2262 = offsetQ_5 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@809.8]
  assign _T_2263 = _T_2261 & _T_2262; // @[AxiStoreQueue.scala 102:61:@810.8]
  assign _T_2266 = io_loadHead <= offsetQ_5; // @[AxiStoreQueue.scala 105:23:@816.10]
  assign _T_2267 = offsetQ_5 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@817.10]
  assign _T_2268 = _T_2266 & _T_2267; // @[AxiStoreQueue.scala 105:49:@818.10]
  assign _T_2270 = _T_2268 == 1'h0; // @[AxiStoreQueue.scala 105:9:@819.10]
  assign _T_2271 = _T_2115 & _T_2270; // @[AxiStoreQueue.scala 104:49:@820.10]
  assign _GEN_660 = _T_2271 ? 1'h0 : checkBits_5; // @[AxiStoreQueue.scala 105:96:@821.10]
  assign _GEN_661 = _T_2263 ? 1'h0 : _GEN_660; // @[AxiStoreQueue.scala 102:102:@811.8]
  assign _GEN_662 = io_loadEmpty ? 1'h0 : _GEN_661; // @[AxiStoreQueue.scala 100:26:@804.6]
  assign _GEN_663 = initBits_5 ? _T_2259 : _GEN_662; // @[AxiStoreQueue.scala 96:35:@789.4]
  assign _T_2284 = _GEN_219 + 4'h1; // @[util.scala 10:8:@832.6]
  assign _GEN_54 = _T_2284 % 5'h10; // @[util.scala 10:14:@833.6]
  assign _T_2285 = _GEN_54[4:0]; // @[util.scala 10:14:@833.6]
  assign _T_2286 = _T_2285 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@834.6]
  assign _T_2287 = io_loadEmpty & _T_2286; // @[AxiStoreQueue.scala 97:50:@835.6]
  assign _T_2289 = _T_2287 == 1'h0; // @[AxiStoreQueue.scala 97:35:@836.6]
  assign _T_2291 = previousLoadHead <= offsetQ_6; // @[AxiStoreQueue.scala 102:35:@844.8]
  assign _T_2292 = offsetQ_6 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@845.8]
  assign _T_2293 = _T_2291 & _T_2292; // @[AxiStoreQueue.scala 102:61:@846.8]
  assign _T_2296 = io_loadHead <= offsetQ_6; // @[AxiStoreQueue.scala 105:23:@852.10]
  assign _T_2297 = offsetQ_6 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@853.10]
  assign _T_2298 = _T_2296 & _T_2297; // @[AxiStoreQueue.scala 105:49:@854.10]
  assign _T_2300 = _T_2298 == 1'h0; // @[AxiStoreQueue.scala 105:9:@855.10]
  assign _T_2301 = _T_2115 & _T_2300; // @[AxiStoreQueue.scala 104:49:@856.10]
  assign _GEN_680 = _T_2301 ? 1'h0 : checkBits_6; // @[AxiStoreQueue.scala 105:96:@857.10]
  assign _GEN_681 = _T_2293 ? 1'h0 : _GEN_680; // @[AxiStoreQueue.scala 102:102:@847.8]
  assign _GEN_682 = io_loadEmpty ? 1'h0 : _GEN_681; // @[AxiStoreQueue.scala 100:26:@840.6]
  assign _GEN_683 = initBits_6 ? _T_2289 : _GEN_682; // @[AxiStoreQueue.scala 96:35:@825.4]
  assign _T_2314 = _GEN_253 + 4'h1; // @[util.scala 10:8:@868.6]
  assign _GEN_55 = _T_2314 % 5'h10; // @[util.scala 10:14:@869.6]
  assign _T_2315 = _GEN_55[4:0]; // @[util.scala 10:14:@869.6]
  assign _T_2316 = _T_2315 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@870.6]
  assign _T_2317 = io_loadEmpty & _T_2316; // @[AxiStoreQueue.scala 97:50:@871.6]
  assign _T_2319 = _T_2317 == 1'h0; // @[AxiStoreQueue.scala 97:35:@872.6]
  assign _T_2321 = previousLoadHead <= offsetQ_7; // @[AxiStoreQueue.scala 102:35:@880.8]
  assign _T_2322 = offsetQ_7 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@881.8]
  assign _T_2323 = _T_2321 & _T_2322; // @[AxiStoreQueue.scala 102:61:@882.8]
  assign _T_2326 = io_loadHead <= offsetQ_7; // @[AxiStoreQueue.scala 105:23:@888.10]
  assign _T_2327 = offsetQ_7 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@889.10]
  assign _T_2328 = _T_2326 & _T_2327; // @[AxiStoreQueue.scala 105:49:@890.10]
  assign _T_2330 = _T_2328 == 1'h0; // @[AxiStoreQueue.scala 105:9:@891.10]
  assign _T_2331 = _T_2115 & _T_2330; // @[AxiStoreQueue.scala 104:49:@892.10]
  assign _GEN_700 = _T_2331 ? 1'h0 : checkBits_7; // @[AxiStoreQueue.scala 105:96:@893.10]
  assign _GEN_701 = _T_2323 ? 1'h0 : _GEN_700; // @[AxiStoreQueue.scala 102:102:@883.8]
  assign _GEN_702 = io_loadEmpty ? 1'h0 : _GEN_701; // @[AxiStoreQueue.scala 100:26:@876.6]
  assign _GEN_703 = initBits_7 ? _T_2319 : _GEN_702; // @[AxiStoreQueue.scala 96:35:@861.4]
  assign _T_2344 = _GEN_287 + 4'h1; // @[util.scala 10:8:@904.6]
  assign _GEN_56 = _T_2344 % 5'h10; // @[util.scala 10:14:@905.6]
  assign _T_2345 = _GEN_56[4:0]; // @[util.scala 10:14:@905.6]
  assign _T_2346 = _T_2345 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@906.6]
  assign _T_2347 = io_loadEmpty & _T_2346; // @[AxiStoreQueue.scala 97:50:@907.6]
  assign _T_2349 = _T_2347 == 1'h0; // @[AxiStoreQueue.scala 97:35:@908.6]
  assign _T_2351 = previousLoadHead <= offsetQ_8; // @[AxiStoreQueue.scala 102:35:@916.8]
  assign _T_2352 = offsetQ_8 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@917.8]
  assign _T_2353 = _T_2351 & _T_2352; // @[AxiStoreQueue.scala 102:61:@918.8]
  assign _T_2356 = io_loadHead <= offsetQ_8; // @[AxiStoreQueue.scala 105:23:@924.10]
  assign _T_2357 = offsetQ_8 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@925.10]
  assign _T_2358 = _T_2356 & _T_2357; // @[AxiStoreQueue.scala 105:49:@926.10]
  assign _T_2360 = _T_2358 == 1'h0; // @[AxiStoreQueue.scala 105:9:@927.10]
  assign _T_2361 = _T_2115 & _T_2360; // @[AxiStoreQueue.scala 104:49:@928.10]
  assign _GEN_720 = _T_2361 ? 1'h0 : checkBits_8; // @[AxiStoreQueue.scala 105:96:@929.10]
  assign _GEN_721 = _T_2353 ? 1'h0 : _GEN_720; // @[AxiStoreQueue.scala 102:102:@919.8]
  assign _GEN_722 = io_loadEmpty ? 1'h0 : _GEN_721; // @[AxiStoreQueue.scala 100:26:@912.6]
  assign _GEN_723 = initBits_8 ? _T_2349 : _GEN_722; // @[AxiStoreQueue.scala 96:35:@897.4]
  assign _T_2374 = _GEN_321 + 4'h1; // @[util.scala 10:8:@940.6]
  assign _GEN_57 = _T_2374 % 5'h10; // @[util.scala 10:14:@941.6]
  assign _T_2375 = _GEN_57[4:0]; // @[util.scala 10:14:@941.6]
  assign _T_2376 = _T_2375 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@942.6]
  assign _T_2377 = io_loadEmpty & _T_2376; // @[AxiStoreQueue.scala 97:50:@943.6]
  assign _T_2379 = _T_2377 == 1'h0; // @[AxiStoreQueue.scala 97:35:@944.6]
  assign _T_2381 = previousLoadHead <= offsetQ_9; // @[AxiStoreQueue.scala 102:35:@952.8]
  assign _T_2382 = offsetQ_9 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@953.8]
  assign _T_2383 = _T_2381 & _T_2382; // @[AxiStoreQueue.scala 102:61:@954.8]
  assign _T_2386 = io_loadHead <= offsetQ_9; // @[AxiStoreQueue.scala 105:23:@960.10]
  assign _T_2387 = offsetQ_9 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@961.10]
  assign _T_2388 = _T_2386 & _T_2387; // @[AxiStoreQueue.scala 105:49:@962.10]
  assign _T_2390 = _T_2388 == 1'h0; // @[AxiStoreQueue.scala 105:9:@963.10]
  assign _T_2391 = _T_2115 & _T_2390; // @[AxiStoreQueue.scala 104:49:@964.10]
  assign _GEN_740 = _T_2391 ? 1'h0 : checkBits_9; // @[AxiStoreQueue.scala 105:96:@965.10]
  assign _GEN_741 = _T_2383 ? 1'h0 : _GEN_740; // @[AxiStoreQueue.scala 102:102:@955.8]
  assign _GEN_742 = io_loadEmpty ? 1'h0 : _GEN_741; // @[AxiStoreQueue.scala 100:26:@948.6]
  assign _GEN_743 = initBits_9 ? _T_2379 : _GEN_742; // @[AxiStoreQueue.scala 96:35:@933.4]
  assign _T_2404 = _GEN_355 + 4'h1; // @[util.scala 10:8:@976.6]
  assign _GEN_58 = _T_2404 % 5'h10; // @[util.scala 10:14:@977.6]
  assign _T_2405 = _GEN_58[4:0]; // @[util.scala 10:14:@977.6]
  assign _T_2406 = _T_2405 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@978.6]
  assign _T_2407 = io_loadEmpty & _T_2406; // @[AxiStoreQueue.scala 97:50:@979.6]
  assign _T_2409 = _T_2407 == 1'h0; // @[AxiStoreQueue.scala 97:35:@980.6]
  assign _T_2411 = previousLoadHead <= offsetQ_10; // @[AxiStoreQueue.scala 102:35:@988.8]
  assign _T_2412 = offsetQ_10 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@989.8]
  assign _T_2413 = _T_2411 & _T_2412; // @[AxiStoreQueue.scala 102:61:@990.8]
  assign _T_2416 = io_loadHead <= offsetQ_10; // @[AxiStoreQueue.scala 105:23:@996.10]
  assign _T_2417 = offsetQ_10 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@997.10]
  assign _T_2418 = _T_2416 & _T_2417; // @[AxiStoreQueue.scala 105:49:@998.10]
  assign _T_2420 = _T_2418 == 1'h0; // @[AxiStoreQueue.scala 105:9:@999.10]
  assign _T_2421 = _T_2115 & _T_2420; // @[AxiStoreQueue.scala 104:49:@1000.10]
  assign _GEN_760 = _T_2421 ? 1'h0 : checkBits_10; // @[AxiStoreQueue.scala 105:96:@1001.10]
  assign _GEN_761 = _T_2413 ? 1'h0 : _GEN_760; // @[AxiStoreQueue.scala 102:102:@991.8]
  assign _GEN_762 = io_loadEmpty ? 1'h0 : _GEN_761; // @[AxiStoreQueue.scala 100:26:@984.6]
  assign _GEN_763 = initBits_10 ? _T_2409 : _GEN_762; // @[AxiStoreQueue.scala 96:35:@969.4]
  assign _T_2434 = _GEN_389 + 4'h1; // @[util.scala 10:8:@1012.6]
  assign _GEN_59 = _T_2434 % 5'h10; // @[util.scala 10:14:@1013.6]
  assign _T_2435 = _GEN_59[4:0]; // @[util.scala 10:14:@1013.6]
  assign _T_2436 = _T_2435 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@1014.6]
  assign _T_2437 = io_loadEmpty & _T_2436; // @[AxiStoreQueue.scala 97:50:@1015.6]
  assign _T_2439 = _T_2437 == 1'h0; // @[AxiStoreQueue.scala 97:35:@1016.6]
  assign _T_2441 = previousLoadHead <= offsetQ_11; // @[AxiStoreQueue.scala 102:35:@1024.8]
  assign _T_2442 = offsetQ_11 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@1025.8]
  assign _T_2443 = _T_2441 & _T_2442; // @[AxiStoreQueue.scala 102:61:@1026.8]
  assign _T_2446 = io_loadHead <= offsetQ_11; // @[AxiStoreQueue.scala 105:23:@1032.10]
  assign _T_2447 = offsetQ_11 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@1033.10]
  assign _T_2448 = _T_2446 & _T_2447; // @[AxiStoreQueue.scala 105:49:@1034.10]
  assign _T_2450 = _T_2448 == 1'h0; // @[AxiStoreQueue.scala 105:9:@1035.10]
  assign _T_2451 = _T_2115 & _T_2450; // @[AxiStoreQueue.scala 104:49:@1036.10]
  assign _GEN_780 = _T_2451 ? 1'h0 : checkBits_11; // @[AxiStoreQueue.scala 105:96:@1037.10]
  assign _GEN_781 = _T_2443 ? 1'h0 : _GEN_780; // @[AxiStoreQueue.scala 102:102:@1027.8]
  assign _GEN_782 = io_loadEmpty ? 1'h0 : _GEN_781; // @[AxiStoreQueue.scala 100:26:@1020.6]
  assign _GEN_783 = initBits_11 ? _T_2439 : _GEN_782; // @[AxiStoreQueue.scala 96:35:@1005.4]
  assign _T_2464 = _GEN_423 + 4'h1; // @[util.scala 10:8:@1048.6]
  assign _GEN_60 = _T_2464 % 5'h10; // @[util.scala 10:14:@1049.6]
  assign _T_2465 = _GEN_60[4:0]; // @[util.scala 10:14:@1049.6]
  assign _T_2466 = _T_2465 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@1050.6]
  assign _T_2467 = io_loadEmpty & _T_2466; // @[AxiStoreQueue.scala 97:50:@1051.6]
  assign _T_2469 = _T_2467 == 1'h0; // @[AxiStoreQueue.scala 97:35:@1052.6]
  assign _T_2471 = previousLoadHead <= offsetQ_12; // @[AxiStoreQueue.scala 102:35:@1060.8]
  assign _T_2472 = offsetQ_12 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@1061.8]
  assign _T_2473 = _T_2471 & _T_2472; // @[AxiStoreQueue.scala 102:61:@1062.8]
  assign _T_2476 = io_loadHead <= offsetQ_12; // @[AxiStoreQueue.scala 105:23:@1068.10]
  assign _T_2477 = offsetQ_12 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@1069.10]
  assign _T_2478 = _T_2476 & _T_2477; // @[AxiStoreQueue.scala 105:49:@1070.10]
  assign _T_2480 = _T_2478 == 1'h0; // @[AxiStoreQueue.scala 105:9:@1071.10]
  assign _T_2481 = _T_2115 & _T_2480; // @[AxiStoreQueue.scala 104:49:@1072.10]
  assign _GEN_800 = _T_2481 ? 1'h0 : checkBits_12; // @[AxiStoreQueue.scala 105:96:@1073.10]
  assign _GEN_801 = _T_2473 ? 1'h0 : _GEN_800; // @[AxiStoreQueue.scala 102:102:@1063.8]
  assign _GEN_802 = io_loadEmpty ? 1'h0 : _GEN_801; // @[AxiStoreQueue.scala 100:26:@1056.6]
  assign _GEN_803 = initBits_12 ? _T_2469 : _GEN_802; // @[AxiStoreQueue.scala 96:35:@1041.4]
  assign _T_2494 = _GEN_457 + 4'h1; // @[util.scala 10:8:@1084.6]
  assign _GEN_61 = _T_2494 % 5'h10; // @[util.scala 10:14:@1085.6]
  assign _T_2495 = _GEN_61[4:0]; // @[util.scala 10:14:@1085.6]
  assign _T_2496 = _T_2495 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@1086.6]
  assign _T_2497 = io_loadEmpty & _T_2496; // @[AxiStoreQueue.scala 97:50:@1087.6]
  assign _T_2499 = _T_2497 == 1'h0; // @[AxiStoreQueue.scala 97:35:@1088.6]
  assign _T_2501 = previousLoadHead <= offsetQ_13; // @[AxiStoreQueue.scala 102:35:@1096.8]
  assign _T_2502 = offsetQ_13 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@1097.8]
  assign _T_2503 = _T_2501 & _T_2502; // @[AxiStoreQueue.scala 102:61:@1098.8]
  assign _T_2506 = io_loadHead <= offsetQ_13; // @[AxiStoreQueue.scala 105:23:@1104.10]
  assign _T_2507 = offsetQ_13 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@1105.10]
  assign _T_2508 = _T_2506 & _T_2507; // @[AxiStoreQueue.scala 105:49:@1106.10]
  assign _T_2510 = _T_2508 == 1'h0; // @[AxiStoreQueue.scala 105:9:@1107.10]
  assign _T_2511 = _T_2115 & _T_2510; // @[AxiStoreQueue.scala 104:49:@1108.10]
  assign _GEN_820 = _T_2511 ? 1'h0 : checkBits_13; // @[AxiStoreQueue.scala 105:96:@1109.10]
  assign _GEN_821 = _T_2503 ? 1'h0 : _GEN_820; // @[AxiStoreQueue.scala 102:102:@1099.8]
  assign _GEN_822 = io_loadEmpty ? 1'h0 : _GEN_821; // @[AxiStoreQueue.scala 100:26:@1092.6]
  assign _GEN_823 = initBits_13 ? _T_2499 : _GEN_822; // @[AxiStoreQueue.scala 96:35:@1077.4]
  assign _T_2524 = _GEN_491 + 4'h1; // @[util.scala 10:8:@1120.6]
  assign _GEN_62 = _T_2524 % 5'h10; // @[util.scala 10:14:@1121.6]
  assign _T_2525 = _GEN_62[4:0]; // @[util.scala 10:14:@1121.6]
  assign _T_2526 = _T_2525 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@1122.6]
  assign _T_2527 = io_loadEmpty & _T_2526; // @[AxiStoreQueue.scala 97:50:@1123.6]
  assign _T_2529 = _T_2527 == 1'h0; // @[AxiStoreQueue.scala 97:35:@1124.6]
  assign _T_2531 = previousLoadHead <= offsetQ_14; // @[AxiStoreQueue.scala 102:35:@1132.8]
  assign _T_2532 = offsetQ_14 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@1133.8]
  assign _T_2533 = _T_2531 & _T_2532; // @[AxiStoreQueue.scala 102:61:@1134.8]
  assign _T_2536 = io_loadHead <= offsetQ_14; // @[AxiStoreQueue.scala 105:23:@1140.10]
  assign _T_2537 = offsetQ_14 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@1141.10]
  assign _T_2538 = _T_2536 & _T_2537; // @[AxiStoreQueue.scala 105:49:@1142.10]
  assign _T_2540 = _T_2538 == 1'h0; // @[AxiStoreQueue.scala 105:9:@1143.10]
  assign _T_2541 = _T_2115 & _T_2540; // @[AxiStoreQueue.scala 104:49:@1144.10]
  assign _GEN_840 = _T_2541 ? 1'h0 : checkBits_14; // @[AxiStoreQueue.scala 105:96:@1145.10]
  assign _GEN_841 = _T_2533 ? 1'h0 : _GEN_840; // @[AxiStoreQueue.scala 102:102:@1135.8]
  assign _GEN_842 = io_loadEmpty ? 1'h0 : _GEN_841; // @[AxiStoreQueue.scala 100:26:@1128.6]
  assign _GEN_843 = initBits_14 ? _T_2529 : _GEN_842; // @[AxiStoreQueue.scala 96:35:@1113.4]
  assign _T_2554 = _GEN_525 + 4'h1; // @[util.scala 10:8:@1156.6]
  assign _GEN_63 = _T_2554 % 5'h10; // @[util.scala 10:14:@1157.6]
  assign _T_2555 = _GEN_63[4:0]; // @[util.scala 10:14:@1157.6]
  assign _T_2556 = _T_2555 == _GEN_1220; // @[AxiStoreQueue.scala 98:56:@1158.6]
  assign _T_2557 = io_loadEmpty & _T_2556; // @[AxiStoreQueue.scala 97:50:@1159.6]
  assign _T_2559 = _T_2557 == 1'h0; // @[AxiStoreQueue.scala 97:35:@1160.6]
  assign _T_2561 = previousLoadHead <= offsetQ_15; // @[AxiStoreQueue.scala 102:35:@1168.8]
  assign _T_2562 = offsetQ_15 < io_loadHead; // @[AxiStoreQueue.scala 102:87:@1169.8]
  assign _T_2563 = _T_2561 & _T_2562; // @[AxiStoreQueue.scala 102:61:@1170.8]
  assign _T_2566 = io_loadHead <= offsetQ_15; // @[AxiStoreQueue.scala 105:23:@1176.10]
  assign _T_2567 = offsetQ_15 < previousLoadHead; // @[AxiStoreQueue.scala 105:75:@1177.10]
  assign _T_2568 = _T_2566 & _T_2567; // @[AxiStoreQueue.scala 105:49:@1178.10]
  assign _T_2570 = _T_2568 == 1'h0; // @[AxiStoreQueue.scala 105:9:@1179.10]
  assign _T_2571 = _T_2115 & _T_2570; // @[AxiStoreQueue.scala 104:49:@1180.10]
  assign _GEN_860 = _T_2571 ? 1'h0 : checkBits_15; // @[AxiStoreQueue.scala 105:96:@1181.10]
  assign _GEN_861 = _T_2563 ? 1'h0 : _GEN_860; // @[AxiStoreQueue.scala 102:102:@1171.8]
  assign _GEN_862 = io_loadEmpty ? 1'h0 : _GEN_861; // @[AxiStoreQueue.scala 100:26:@1164.6]
  assign _GEN_863 = initBits_15 ? _T_2559 : _GEN_862; // @[AxiStoreQueue.scala 96:35:@1149.4]
  assign _T_2573 = io_loadHead < io_loadTail; // @[AxiStoreQueue.scala 121:103:@1185.4]
  assign _T_2575 = io_loadHead <= 4'h0; // @[AxiStoreQueue.scala 122:17:@1186.4]
  assign _T_2577 = 4'h0 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1187.4]
  assign _T_2578 = _T_2575 & _T_2577; // @[AxiStoreQueue.scala 122:26:@1188.4]
  assign _T_2580 = io_loadEmpty == 1'h0; // @[AxiStoreQueue.scala 122:50:@1189.4]
  assign _T_2582 = io_loadTail <= 4'h0; // @[AxiStoreQueue.scala 122:81:@1190.4]
  assign _T_2584 = 4'h0 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1191.4]
  assign _T_2585 = _T_2582 & _T_2584; // @[AxiStoreQueue.scala 122:90:@1192.4]
  assign _T_2587 = _T_2585 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1193.4]
  assign _T_2588 = _T_2580 & _T_2587; // @[AxiStoreQueue.scala 122:64:@1194.4]
  assign validEntriesInLoadQ_0 = _T_2573 ? _T_2578 : _T_2588; // @[AxiStoreQueue.scala 121:90:@1195.4]
  assign _T_2592 = io_loadHead <= 4'h1; // @[AxiStoreQueue.scala 122:17:@1197.4]
  assign _T_2594 = 4'h1 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1198.4]
  assign _T_2595 = _T_2592 & _T_2594; // @[AxiStoreQueue.scala 122:26:@1199.4]
  assign _T_2599 = io_loadTail <= 4'h1; // @[AxiStoreQueue.scala 122:81:@1201.4]
  assign _T_2601 = 4'h1 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1202.4]
  assign _T_2602 = _T_2599 & _T_2601; // @[AxiStoreQueue.scala 122:90:@1203.4]
  assign _T_2604 = _T_2602 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1204.4]
  assign _T_2605 = _T_2580 & _T_2604; // @[AxiStoreQueue.scala 122:64:@1205.4]
  assign validEntriesInLoadQ_1 = _T_2573 ? _T_2595 : _T_2605; // @[AxiStoreQueue.scala 121:90:@1206.4]
  assign _T_2609 = io_loadHead <= 4'h2; // @[AxiStoreQueue.scala 122:17:@1208.4]
  assign _T_2611 = 4'h2 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1209.4]
  assign _T_2612 = _T_2609 & _T_2611; // @[AxiStoreQueue.scala 122:26:@1210.4]
  assign _T_2616 = io_loadTail <= 4'h2; // @[AxiStoreQueue.scala 122:81:@1212.4]
  assign _T_2618 = 4'h2 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1213.4]
  assign _T_2619 = _T_2616 & _T_2618; // @[AxiStoreQueue.scala 122:90:@1214.4]
  assign _T_2621 = _T_2619 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1215.4]
  assign _T_2622 = _T_2580 & _T_2621; // @[AxiStoreQueue.scala 122:64:@1216.4]
  assign validEntriesInLoadQ_2 = _T_2573 ? _T_2612 : _T_2622; // @[AxiStoreQueue.scala 121:90:@1217.4]
  assign _T_2626 = io_loadHead <= 4'h3; // @[AxiStoreQueue.scala 122:17:@1219.4]
  assign _T_2628 = 4'h3 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1220.4]
  assign _T_2629 = _T_2626 & _T_2628; // @[AxiStoreQueue.scala 122:26:@1221.4]
  assign _T_2633 = io_loadTail <= 4'h3; // @[AxiStoreQueue.scala 122:81:@1223.4]
  assign _T_2635 = 4'h3 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1224.4]
  assign _T_2636 = _T_2633 & _T_2635; // @[AxiStoreQueue.scala 122:90:@1225.4]
  assign _T_2638 = _T_2636 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1226.4]
  assign _T_2639 = _T_2580 & _T_2638; // @[AxiStoreQueue.scala 122:64:@1227.4]
  assign validEntriesInLoadQ_3 = _T_2573 ? _T_2629 : _T_2639; // @[AxiStoreQueue.scala 121:90:@1228.4]
  assign _T_2643 = io_loadHead <= 4'h4; // @[AxiStoreQueue.scala 122:17:@1230.4]
  assign _T_2645 = 4'h4 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1231.4]
  assign _T_2646 = _T_2643 & _T_2645; // @[AxiStoreQueue.scala 122:26:@1232.4]
  assign _T_2650 = io_loadTail <= 4'h4; // @[AxiStoreQueue.scala 122:81:@1234.4]
  assign _T_2652 = 4'h4 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1235.4]
  assign _T_2653 = _T_2650 & _T_2652; // @[AxiStoreQueue.scala 122:90:@1236.4]
  assign _T_2655 = _T_2653 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1237.4]
  assign _T_2656 = _T_2580 & _T_2655; // @[AxiStoreQueue.scala 122:64:@1238.4]
  assign validEntriesInLoadQ_4 = _T_2573 ? _T_2646 : _T_2656; // @[AxiStoreQueue.scala 121:90:@1239.4]
  assign _T_2660 = io_loadHead <= 4'h5; // @[AxiStoreQueue.scala 122:17:@1241.4]
  assign _T_2662 = 4'h5 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1242.4]
  assign _T_2663 = _T_2660 & _T_2662; // @[AxiStoreQueue.scala 122:26:@1243.4]
  assign _T_2667 = io_loadTail <= 4'h5; // @[AxiStoreQueue.scala 122:81:@1245.4]
  assign _T_2669 = 4'h5 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1246.4]
  assign _T_2670 = _T_2667 & _T_2669; // @[AxiStoreQueue.scala 122:90:@1247.4]
  assign _T_2672 = _T_2670 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1248.4]
  assign _T_2673 = _T_2580 & _T_2672; // @[AxiStoreQueue.scala 122:64:@1249.4]
  assign validEntriesInLoadQ_5 = _T_2573 ? _T_2663 : _T_2673; // @[AxiStoreQueue.scala 121:90:@1250.4]
  assign _T_2677 = io_loadHead <= 4'h6; // @[AxiStoreQueue.scala 122:17:@1252.4]
  assign _T_2679 = 4'h6 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1253.4]
  assign _T_2680 = _T_2677 & _T_2679; // @[AxiStoreQueue.scala 122:26:@1254.4]
  assign _T_2684 = io_loadTail <= 4'h6; // @[AxiStoreQueue.scala 122:81:@1256.4]
  assign _T_2686 = 4'h6 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1257.4]
  assign _T_2687 = _T_2684 & _T_2686; // @[AxiStoreQueue.scala 122:90:@1258.4]
  assign _T_2689 = _T_2687 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1259.4]
  assign _T_2690 = _T_2580 & _T_2689; // @[AxiStoreQueue.scala 122:64:@1260.4]
  assign validEntriesInLoadQ_6 = _T_2573 ? _T_2680 : _T_2690; // @[AxiStoreQueue.scala 121:90:@1261.4]
  assign _T_2694 = io_loadHead <= 4'h7; // @[AxiStoreQueue.scala 122:17:@1263.4]
  assign _T_2696 = 4'h7 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1264.4]
  assign _T_2697 = _T_2694 & _T_2696; // @[AxiStoreQueue.scala 122:26:@1265.4]
  assign _T_2701 = io_loadTail <= 4'h7; // @[AxiStoreQueue.scala 122:81:@1267.4]
  assign _T_2703 = 4'h7 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1268.4]
  assign _T_2704 = _T_2701 & _T_2703; // @[AxiStoreQueue.scala 122:90:@1269.4]
  assign _T_2706 = _T_2704 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1270.4]
  assign _T_2707 = _T_2580 & _T_2706; // @[AxiStoreQueue.scala 122:64:@1271.4]
  assign validEntriesInLoadQ_7 = _T_2573 ? _T_2697 : _T_2707; // @[AxiStoreQueue.scala 121:90:@1272.4]
  assign _T_2711 = io_loadHead <= 4'h8; // @[AxiStoreQueue.scala 122:17:@1274.4]
  assign _T_2713 = 4'h8 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1275.4]
  assign _T_2714 = _T_2711 & _T_2713; // @[AxiStoreQueue.scala 122:26:@1276.4]
  assign _T_2718 = io_loadTail <= 4'h8; // @[AxiStoreQueue.scala 122:81:@1278.4]
  assign _T_2720 = 4'h8 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1279.4]
  assign _T_2721 = _T_2718 & _T_2720; // @[AxiStoreQueue.scala 122:90:@1280.4]
  assign _T_2723 = _T_2721 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1281.4]
  assign _T_2724 = _T_2580 & _T_2723; // @[AxiStoreQueue.scala 122:64:@1282.4]
  assign validEntriesInLoadQ_8 = _T_2573 ? _T_2714 : _T_2724; // @[AxiStoreQueue.scala 121:90:@1283.4]
  assign _T_2728 = io_loadHead <= 4'h9; // @[AxiStoreQueue.scala 122:17:@1285.4]
  assign _T_2730 = 4'h9 < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1286.4]
  assign _T_2731 = _T_2728 & _T_2730; // @[AxiStoreQueue.scala 122:26:@1287.4]
  assign _T_2735 = io_loadTail <= 4'h9; // @[AxiStoreQueue.scala 122:81:@1289.4]
  assign _T_2737 = 4'h9 < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1290.4]
  assign _T_2738 = _T_2735 & _T_2737; // @[AxiStoreQueue.scala 122:90:@1291.4]
  assign _T_2740 = _T_2738 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1292.4]
  assign _T_2741 = _T_2580 & _T_2740; // @[AxiStoreQueue.scala 122:64:@1293.4]
  assign validEntriesInLoadQ_9 = _T_2573 ? _T_2731 : _T_2741; // @[AxiStoreQueue.scala 121:90:@1294.4]
  assign _T_2745 = io_loadHead <= 4'ha; // @[AxiStoreQueue.scala 122:17:@1296.4]
  assign _T_2747 = 4'ha < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1297.4]
  assign _T_2748 = _T_2745 & _T_2747; // @[AxiStoreQueue.scala 122:26:@1298.4]
  assign _T_2752 = io_loadTail <= 4'ha; // @[AxiStoreQueue.scala 122:81:@1300.4]
  assign _T_2754 = 4'ha < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1301.4]
  assign _T_2755 = _T_2752 & _T_2754; // @[AxiStoreQueue.scala 122:90:@1302.4]
  assign _T_2757 = _T_2755 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1303.4]
  assign _T_2758 = _T_2580 & _T_2757; // @[AxiStoreQueue.scala 122:64:@1304.4]
  assign validEntriesInLoadQ_10 = _T_2573 ? _T_2748 : _T_2758; // @[AxiStoreQueue.scala 121:90:@1305.4]
  assign _T_2762 = io_loadHead <= 4'hb; // @[AxiStoreQueue.scala 122:17:@1307.4]
  assign _T_2764 = 4'hb < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1308.4]
  assign _T_2765 = _T_2762 & _T_2764; // @[AxiStoreQueue.scala 122:26:@1309.4]
  assign _T_2769 = io_loadTail <= 4'hb; // @[AxiStoreQueue.scala 122:81:@1311.4]
  assign _T_2771 = 4'hb < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1312.4]
  assign _T_2772 = _T_2769 & _T_2771; // @[AxiStoreQueue.scala 122:90:@1313.4]
  assign _T_2774 = _T_2772 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1314.4]
  assign _T_2775 = _T_2580 & _T_2774; // @[AxiStoreQueue.scala 122:64:@1315.4]
  assign validEntriesInLoadQ_11 = _T_2573 ? _T_2765 : _T_2775; // @[AxiStoreQueue.scala 121:90:@1316.4]
  assign _T_2779 = io_loadHead <= 4'hc; // @[AxiStoreQueue.scala 122:17:@1318.4]
  assign _T_2781 = 4'hc < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1319.4]
  assign _T_2782 = _T_2779 & _T_2781; // @[AxiStoreQueue.scala 122:26:@1320.4]
  assign _T_2786 = io_loadTail <= 4'hc; // @[AxiStoreQueue.scala 122:81:@1322.4]
  assign _T_2788 = 4'hc < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1323.4]
  assign _T_2789 = _T_2786 & _T_2788; // @[AxiStoreQueue.scala 122:90:@1324.4]
  assign _T_2791 = _T_2789 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1325.4]
  assign _T_2792 = _T_2580 & _T_2791; // @[AxiStoreQueue.scala 122:64:@1326.4]
  assign validEntriesInLoadQ_12 = _T_2573 ? _T_2782 : _T_2792; // @[AxiStoreQueue.scala 121:90:@1327.4]
  assign _T_2796 = io_loadHead <= 4'hd; // @[AxiStoreQueue.scala 122:17:@1329.4]
  assign _T_2798 = 4'hd < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1330.4]
  assign _T_2799 = _T_2796 & _T_2798; // @[AxiStoreQueue.scala 122:26:@1331.4]
  assign _T_2803 = io_loadTail <= 4'hd; // @[AxiStoreQueue.scala 122:81:@1333.4]
  assign _T_2805 = 4'hd < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1334.4]
  assign _T_2806 = _T_2803 & _T_2805; // @[AxiStoreQueue.scala 122:90:@1335.4]
  assign _T_2808 = _T_2806 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1336.4]
  assign _T_2809 = _T_2580 & _T_2808; // @[AxiStoreQueue.scala 122:64:@1337.4]
  assign validEntriesInLoadQ_13 = _T_2573 ? _T_2799 : _T_2809; // @[AxiStoreQueue.scala 121:90:@1338.4]
  assign _T_2813 = io_loadHead <= 4'he; // @[AxiStoreQueue.scala 122:17:@1340.4]
  assign _T_2815 = 4'he < io_loadTail; // @[AxiStoreQueue.scala 122:35:@1341.4]
  assign _T_2816 = _T_2813 & _T_2815; // @[AxiStoreQueue.scala 122:26:@1342.4]
  assign _T_2820 = io_loadTail <= 4'he; // @[AxiStoreQueue.scala 122:81:@1344.4]
  assign _T_2822 = 4'he < io_loadHead; // @[AxiStoreQueue.scala 122:99:@1345.4]
  assign _T_2823 = _T_2820 & _T_2822; // @[AxiStoreQueue.scala 122:90:@1346.4]
  assign _T_2825 = _T_2823 == 1'h0; // @[AxiStoreQueue.scala 122:67:@1347.4]
  assign _T_2826 = _T_2580 & _T_2825; // @[AxiStoreQueue.scala 122:64:@1348.4]
  assign validEntriesInLoadQ_14 = _T_2573 ? _T_2816 : _T_2826; // @[AxiStoreQueue.scala 121:90:@1349.4]
  assign validEntriesInLoadQ_15 = _T_2573 ? 1'h0 : _T_2580; // @[AxiStoreQueue.scala 121:90:@1360.4]
  assign _GEN_865 = 4'h1 == dummyHead ? offsetQ_1 : offsetQ_0; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_866 = 4'h2 == dummyHead ? offsetQ_2 : _GEN_865; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_867 = 4'h3 == dummyHead ? offsetQ_3 : _GEN_866; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_868 = 4'h4 == dummyHead ? offsetQ_4 : _GEN_867; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_869 = 4'h5 == dummyHead ? offsetQ_5 : _GEN_868; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_870 = 4'h6 == dummyHead ? offsetQ_6 : _GEN_869; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_871 = 4'h7 == dummyHead ? offsetQ_7 : _GEN_870; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_872 = 4'h8 == dummyHead ? offsetQ_8 : _GEN_871; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_873 = 4'h9 == dummyHead ? offsetQ_9 : _GEN_872; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_874 = 4'ha == dummyHead ? offsetQ_10 : _GEN_873; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_875 = 4'hb == dummyHead ? offsetQ_11 : _GEN_874; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_876 = 4'hc == dummyHead ? offsetQ_12 : _GEN_875; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_877 = 4'hd == dummyHead ? offsetQ_13 : _GEN_876; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_878 = 4'he == dummyHead ? offsetQ_14 : _GEN_877; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _GEN_879 = 4'hf == dummyHead ? offsetQ_15 : _GEN_878; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign _T_2869 = io_loadHead <= _GEN_879; // @[AxiStoreQueue.scala 128:96:@1378.4]
  assign loadsToCheck_0 = _T_2869 ? _T_2575 : 1'h1; // @[AxiStoreQueue.scala 128:83:@1386.4]
  assign _T_2899 = 4'h1 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1389.4]
  assign _T_2900 = _T_2592 & _T_2899; // @[AxiStoreQueue.scala 129:26:@1390.4]
  assign _T_2905 = _GEN_879 < 4'h1; // @[AxiStoreQueue.scala 129:79:@1391.4]
  assign _T_2908 = _T_2905 & _T_2601; // @[AxiStoreQueue.scala 129:87:@1393.4]
  assign _T_2910 = _T_2908 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1394.4]
  assign loadsToCheck_1 = _T_2869 ? _T_2900 : _T_2910; // @[AxiStoreQueue.scala 128:83:@1395.4]
  assign _T_2922 = 4'h2 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1398.4]
  assign _T_2923 = _T_2609 & _T_2922; // @[AxiStoreQueue.scala 129:26:@1399.4]
  assign _T_2928 = _GEN_879 < 4'h2; // @[AxiStoreQueue.scala 129:79:@1400.4]
  assign _T_2931 = _T_2928 & _T_2618; // @[AxiStoreQueue.scala 129:87:@1402.4]
  assign _T_2933 = _T_2931 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1403.4]
  assign loadsToCheck_2 = _T_2869 ? _T_2923 : _T_2933; // @[AxiStoreQueue.scala 128:83:@1404.4]
  assign _T_2945 = 4'h3 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1407.4]
  assign _T_2946 = _T_2626 & _T_2945; // @[AxiStoreQueue.scala 129:26:@1408.4]
  assign _T_2951 = _GEN_879 < 4'h3; // @[AxiStoreQueue.scala 129:79:@1409.4]
  assign _T_2954 = _T_2951 & _T_2635; // @[AxiStoreQueue.scala 129:87:@1411.4]
  assign _T_2956 = _T_2954 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1412.4]
  assign loadsToCheck_3 = _T_2869 ? _T_2946 : _T_2956; // @[AxiStoreQueue.scala 128:83:@1413.4]
  assign _T_2968 = 4'h4 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1416.4]
  assign _T_2969 = _T_2643 & _T_2968; // @[AxiStoreQueue.scala 129:26:@1417.4]
  assign _T_2974 = _GEN_879 < 4'h4; // @[AxiStoreQueue.scala 129:79:@1418.4]
  assign _T_2977 = _T_2974 & _T_2652; // @[AxiStoreQueue.scala 129:87:@1420.4]
  assign _T_2979 = _T_2977 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1421.4]
  assign loadsToCheck_4 = _T_2869 ? _T_2969 : _T_2979; // @[AxiStoreQueue.scala 128:83:@1422.4]
  assign _T_2991 = 4'h5 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1425.4]
  assign _T_2992 = _T_2660 & _T_2991; // @[AxiStoreQueue.scala 129:26:@1426.4]
  assign _T_2997 = _GEN_879 < 4'h5; // @[AxiStoreQueue.scala 129:79:@1427.4]
  assign _T_3000 = _T_2997 & _T_2669; // @[AxiStoreQueue.scala 129:87:@1429.4]
  assign _T_3002 = _T_3000 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1430.4]
  assign loadsToCheck_5 = _T_2869 ? _T_2992 : _T_3002; // @[AxiStoreQueue.scala 128:83:@1431.4]
  assign _T_3014 = 4'h6 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1434.4]
  assign _T_3015 = _T_2677 & _T_3014; // @[AxiStoreQueue.scala 129:26:@1435.4]
  assign _T_3020 = _GEN_879 < 4'h6; // @[AxiStoreQueue.scala 129:79:@1436.4]
  assign _T_3023 = _T_3020 & _T_2686; // @[AxiStoreQueue.scala 129:87:@1438.4]
  assign _T_3025 = _T_3023 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1439.4]
  assign loadsToCheck_6 = _T_2869 ? _T_3015 : _T_3025; // @[AxiStoreQueue.scala 128:83:@1440.4]
  assign _T_3037 = 4'h7 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1443.4]
  assign _T_3038 = _T_2694 & _T_3037; // @[AxiStoreQueue.scala 129:26:@1444.4]
  assign _T_3043 = _GEN_879 < 4'h7; // @[AxiStoreQueue.scala 129:79:@1445.4]
  assign _T_3046 = _T_3043 & _T_2703; // @[AxiStoreQueue.scala 129:87:@1447.4]
  assign _T_3048 = _T_3046 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1448.4]
  assign loadsToCheck_7 = _T_2869 ? _T_3038 : _T_3048; // @[AxiStoreQueue.scala 128:83:@1449.4]
  assign _T_3060 = 4'h8 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1452.4]
  assign _T_3061 = _T_2711 & _T_3060; // @[AxiStoreQueue.scala 129:26:@1453.4]
  assign _T_3066 = _GEN_879 < 4'h8; // @[AxiStoreQueue.scala 129:79:@1454.4]
  assign _T_3069 = _T_3066 & _T_2720; // @[AxiStoreQueue.scala 129:87:@1456.4]
  assign _T_3071 = _T_3069 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1457.4]
  assign loadsToCheck_8 = _T_2869 ? _T_3061 : _T_3071; // @[AxiStoreQueue.scala 128:83:@1458.4]
  assign _T_3083 = 4'h9 <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1461.4]
  assign _T_3084 = _T_2728 & _T_3083; // @[AxiStoreQueue.scala 129:26:@1462.4]
  assign _T_3089 = _GEN_879 < 4'h9; // @[AxiStoreQueue.scala 129:79:@1463.4]
  assign _T_3092 = _T_3089 & _T_2737; // @[AxiStoreQueue.scala 129:87:@1465.4]
  assign _T_3094 = _T_3092 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1466.4]
  assign loadsToCheck_9 = _T_2869 ? _T_3084 : _T_3094; // @[AxiStoreQueue.scala 128:83:@1467.4]
  assign _T_3106 = 4'ha <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1470.4]
  assign _T_3107 = _T_2745 & _T_3106; // @[AxiStoreQueue.scala 129:26:@1471.4]
  assign _T_3112 = _GEN_879 < 4'ha; // @[AxiStoreQueue.scala 129:79:@1472.4]
  assign _T_3115 = _T_3112 & _T_2754; // @[AxiStoreQueue.scala 129:87:@1474.4]
  assign _T_3117 = _T_3115 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1475.4]
  assign loadsToCheck_10 = _T_2869 ? _T_3107 : _T_3117; // @[AxiStoreQueue.scala 128:83:@1476.4]
  assign _T_3129 = 4'hb <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1479.4]
  assign _T_3130 = _T_2762 & _T_3129; // @[AxiStoreQueue.scala 129:26:@1480.4]
  assign _T_3135 = _GEN_879 < 4'hb; // @[AxiStoreQueue.scala 129:79:@1481.4]
  assign _T_3138 = _T_3135 & _T_2771; // @[AxiStoreQueue.scala 129:87:@1483.4]
  assign _T_3140 = _T_3138 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1484.4]
  assign loadsToCheck_11 = _T_2869 ? _T_3130 : _T_3140; // @[AxiStoreQueue.scala 128:83:@1485.4]
  assign _T_3152 = 4'hc <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1488.4]
  assign _T_3153 = _T_2779 & _T_3152; // @[AxiStoreQueue.scala 129:26:@1489.4]
  assign _T_3158 = _GEN_879 < 4'hc; // @[AxiStoreQueue.scala 129:79:@1490.4]
  assign _T_3161 = _T_3158 & _T_2788; // @[AxiStoreQueue.scala 129:87:@1492.4]
  assign _T_3163 = _T_3161 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1493.4]
  assign loadsToCheck_12 = _T_2869 ? _T_3153 : _T_3163; // @[AxiStoreQueue.scala 128:83:@1494.4]
  assign _T_3175 = 4'hd <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1497.4]
  assign _T_3176 = _T_2796 & _T_3175; // @[AxiStoreQueue.scala 129:26:@1498.4]
  assign _T_3181 = _GEN_879 < 4'hd; // @[AxiStoreQueue.scala 129:79:@1499.4]
  assign _T_3184 = _T_3181 & _T_2805; // @[AxiStoreQueue.scala 129:87:@1501.4]
  assign _T_3186 = _T_3184 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1502.4]
  assign loadsToCheck_13 = _T_2869 ? _T_3176 : _T_3186; // @[AxiStoreQueue.scala 128:83:@1503.4]
  assign _T_3198 = 4'he <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1506.4]
  assign _T_3199 = _T_2813 & _T_3198; // @[AxiStoreQueue.scala 129:26:@1507.4]
  assign _T_3204 = _GEN_879 < 4'he; // @[AxiStoreQueue.scala 129:79:@1508.4]
  assign _T_3207 = _T_3204 & _T_2822; // @[AxiStoreQueue.scala 129:87:@1510.4]
  assign _T_3209 = _T_3207 == 1'h0; // @[AxiStoreQueue.scala 129:58:@1511.4]
  assign loadsToCheck_14 = _T_2869 ? _T_3199 : _T_3209; // @[AxiStoreQueue.scala 128:83:@1512.4]
  assign _T_3221 = 4'hf <= _GEN_879; // @[AxiStoreQueue.scala 129:35:@1515.4]
  assign loadsToCheck_15 = _T_2869 ? _T_3221 : 1'h1; // @[AxiStoreQueue.scala 128:83:@1521.4]
  assign _T_3255 = loadsToCheck_0 & validEntriesInLoadQ_0; // @[AxiStoreQueue.scala 135:16:@1539.4]
  assign _GEN_881 = 4'h1 == dummyHead ? checkBits_1 : checkBits_0; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_882 = 4'h2 == dummyHead ? checkBits_2 : _GEN_881; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_883 = 4'h3 == dummyHead ? checkBits_3 : _GEN_882; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_884 = 4'h4 == dummyHead ? checkBits_4 : _GEN_883; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_885 = 4'h5 == dummyHead ? checkBits_5 : _GEN_884; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_886 = 4'h6 == dummyHead ? checkBits_6 : _GEN_885; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_887 = 4'h7 == dummyHead ? checkBits_7 : _GEN_886; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_888 = 4'h8 == dummyHead ? checkBits_8 : _GEN_887; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_889 = 4'h9 == dummyHead ? checkBits_9 : _GEN_888; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_890 = 4'ha == dummyHead ? checkBits_10 : _GEN_889; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_891 = 4'hb == dummyHead ? checkBits_11 : _GEN_890; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_892 = 4'hc == dummyHead ? checkBits_12 : _GEN_891; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_893 = 4'hd == dummyHead ? checkBits_13 : _GEN_892; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_894 = 4'he == dummyHead ? checkBits_14 : _GEN_893; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _GEN_895 = 4'hf == dummyHead ? checkBits_15 : _GEN_894; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign entriesToCheck_0 = _T_3255 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1540.4]
  assign _T_3260 = loadsToCheck_1 & validEntriesInLoadQ_1; // @[AxiStoreQueue.scala 135:16:@1541.4]
  assign entriesToCheck_1 = _T_3260 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1542.4]
  assign _T_3265 = loadsToCheck_2 & validEntriesInLoadQ_2; // @[AxiStoreQueue.scala 135:16:@1543.4]
  assign entriesToCheck_2 = _T_3265 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1544.4]
  assign _T_3270 = loadsToCheck_3 & validEntriesInLoadQ_3; // @[AxiStoreQueue.scala 135:16:@1545.4]
  assign entriesToCheck_3 = _T_3270 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1546.4]
  assign _T_3275 = loadsToCheck_4 & validEntriesInLoadQ_4; // @[AxiStoreQueue.scala 135:16:@1547.4]
  assign entriesToCheck_4 = _T_3275 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1548.4]
  assign _T_3280 = loadsToCheck_5 & validEntriesInLoadQ_5; // @[AxiStoreQueue.scala 135:16:@1549.4]
  assign entriesToCheck_5 = _T_3280 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1550.4]
  assign _T_3285 = loadsToCheck_6 & validEntriesInLoadQ_6; // @[AxiStoreQueue.scala 135:16:@1551.4]
  assign entriesToCheck_6 = _T_3285 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1552.4]
  assign _T_3290 = loadsToCheck_7 & validEntriesInLoadQ_7; // @[AxiStoreQueue.scala 135:16:@1553.4]
  assign entriesToCheck_7 = _T_3290 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1554.4]
  assign _T_3295 = loadsToCheck_8 & validEntriesInLoadQ_8; // @[AxiStoreQueue.scala 135:16:@1555.4]
  assign entriesToCheck_8 = _T_3295 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1556.4]
  assign _T_3300 = loadsToCheck_9 & validEntriesInLoadQ_9; // @[AxiStoreQueue.scala 135:16:@1557.4]
  assign entriesToCheck_9 = _T_3300 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1558.4]
  assign _T_3305 = loadsToCheck_10 & validEntriesInLoadQ_10; // @[AxiStoreQueue.scala 135:16:@1559.4]
  assign entriesToCheck_10 = _T_3305 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1560.4]
  assign _T_3310 = loadsToCheck_11 & validEntriesInLoadQ_11; // @[AxiStoreQueue.scala 135:16:@1561.4]
  assign entriesToCheck_11 = _T_3310 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1562.4]
  assign _T_3315 = loadsToCheck_12 & validEntriesInLoadQ_12; // @[AxiStoreQueue.scala 135:16:@1563.4]
  assign entriesToCheck_12 = _T_3315 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1564.4]
  assign _T_3320 = loadsToCheck_13 & validEntriesInLoadQ_13; // @[AxiStoreQueue.scala 135:16:@1565.4]
  assign entriesToCheck_13 = _T_3320 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1566.4]
  assign _T_3325 = loadsToCheck_14 & validEntriesInLoadQ_14; // @[AxiStoreQueue.scala 135:16:@1567.4]
  assign entriesToCheck_14 = _T_3325 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1568.4]
  assign _T_3330 = loadsToCheck_15 & validEntriesInLoadQ_15; // @[AxiStoreQueue.scala 135:16:@1569.4]
  assign entriesToCheck_15 = _T_3330 & _GEN_895; // @[AxiStoreQueue.scala 135:24:@1570.4]
  assign _T_3378 = entriesToCheck_0 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1589.4]
  assign _T_3379 = _T_3378 | io_loadDataDone_0; // @[AxiStoreQueue.scala 142:64:@1590.4]
  assign _GEN_897 = 4'h1 == dummyHead ? addrQ_1 : addrQ_0; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_898 = 4'h2 == dummyHead ? addrQ_2 : _GEN_897; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_899 = 4'h3 == dummyHead ? addrQ_3 : _GEN_898; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_900 = 4'h4 == dummyHead ? addrQ_4 : _GEN_899; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_901 = 4'h5 == dummyHead ? addrQ_5 : _GEN_900; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_902 = 4'h6 == dummyHead ? addrQ_6 : _GEN_901; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_903 = 4'h7 == dummyHead ? addrQ_7 : _GEN_902; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_904 = 4'h8 == dummyHead ? addrQ_8 : _GEN_903; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_905 = 4'h9 == dummyHead ? addrQ_9 : _GEN_904; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_906 = 4'ha == dummyHead ? addrQ_10 : _GEN_905; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_907 = 4'hb == dummyHead ? addrQ_11 : _GEN_906; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_908 = 4'hc == dummyHead ? addrQ_12 : _GEN_907; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_909 = 4'hd == dummyHead ? addrQ_13 : _GEN_908; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_910 = 4'he == dummyHead ? addrQ_14 : _GEN_909; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _GEN_911 = 4'hf == dummyHead ? addrQ_15 : _GEN_910; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _T_3383 = _GEN_911 != io_loadAddressQueue_0; // @[AxiStoreQueue.scala 143:56:@1591.4]
  assign _T_3384 = io_loadAddressDone_0 & _T_3383; // @[AxiStoreQueue.scala 143:36:@1592.4]
  assign noConflicts_0 = _T_3379 | _T_3384; // @[AxiStoreQueue.scala 142:95:@1593.4]
  assign _T_3387 = entriesToCheck_1 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1595.4]
  assign _T_3388 = _T_3387 | io_loadDataDone_1; // @[AxiStoreQueue.scala 142:64:@1596.4]
  assign _T_3392 = _GEN_911 != io_loadAddressQueue_1; // @[AxiStoreQueue.scala 143:56:@1597.4]
  assign _T_3393 = io_loadAddressDone_1 & _T_3392; // @[AxiStoreQueue.scala 143:36:@1598.4]
  assign noConflicts_1 = _T_3388 | _T_3393; // @[AxiStoreQueue.scala 142:95:@1599.4]
  assign _T_3396 = entriesToCheck_2 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1601.4]
  assign _T_3397 = _T_3396 | io_loadDataDone_2; // @[AxiStoreQueue.scala 142:64:@1602.4]
  assign _T_3401 = _GEN_911 != io_loadAddressQueue_2; // @[AxiStoreQueue.scala 143:56:@1603.4]
  assign _T_3402 = io_loadAddressDone_2 & _T_3401; // @[AxiStoreQueue.scala 143:36:@1604.4]
  assign noConflicts_2 = _T_3397 | _T_3402; // @[AxiStoreQueue.scala 142:95:@1605.4]
  assign _T_3405 = entriesToCheck_3 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1607.4]
  assign _T_3406 = _T_3405 | io_loadDataDone_3; // @[AxiStoreQueue.scala 142:64:@1608.4]
  assign _T_3410 = _GEN_911 != io_loadAddressQueue_3; // @[AxiStoreQueue.scala 143:56:@1609.4]
  assign _T_3411 = io_loadAddressDone_3 & _T_3410; // @[AxiStoreQueue.scala 143:36:@1610.4]
  assign noConflicts_3 = _T_3406 | _T_3411; // @[AxiStoreQueue.scala 142:95:@1611.4]
  assign _T_3414 = entriesToCheck_4 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1613.4]
  assign _T_3415 = _T_3414 | io_loadDataDone_4; // @[AxiStoreQueue.scala 142:64:@1614.4]
  assign _T_3419 = _GEN_911 != io_loadAddressQueue_4; // @[AxiStoreQueue.scala 143:56:@1615.4]
  assign _T_3420 = io_loadAddressDone_4 & _T_3419; // @[AxiStoreQueue.scala 143:36:@1616.4]
  assign noConflicts_4 = _T_3415 | _T_3420; // @[AxiStoreQueue.scala 142:95:@1617.4]
  assign _T_3423 = entriesToCheck_5 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1619.4]
  assign _T_3424 = _T_3423 | io_loadDataDone_5; // @[AxiStoreQueue.scala 142:64:@1620.4]
  assign _T_3428 = _GEN_911 != io_loadAddressQueue_5; // @[AxiStoreQueue.scala 143:56:@1621.4]
  assign _T_3429 = io_loadAddressDone_5 & _T_3428; // @[AxiStoreQueue.scala 143:36:@1622.4]
  assign noConflicts_5 = _T_3424 | _T_3429; // @[AxiStoreQueue.scala 142:95:@1623.4]
  assign _T_3432 = entriesToCheck_6 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1625.4]
  assign _T_3433 = _T_3432 | io_loadDataDone_6; // @[AxiStoreQueue.scala 142:64:@1626.4]
  assign _T_3437 = _GEN_911 != io_loadAddressQueue_6; // @[AxiStoreQueue.scala 143:56:@1627.4]
  assign _T_3438 = io_loadAddressDone_6 & _T_3437; // @[AxiStoreQueue.scala 143:36:@1628.4]
  assign noConflicts_6 = _T_3433 | _T_3438; // @[AxiStoreQueue.scala 142:95:@1629.4]
  assign _T_3441 = entriesToCheck_7 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1631.4]
  assign _T_3442 = _T_3441 | io_loadDataDone_7; // @[AxiStoreQueue.scala 142:64:@1632.4]
  assign _T_3446 = _GEN_911 != io_loadAddressQueue_7; // @[AxiStoreQueue.scala 143:56:@1633.4]
  assign _T_3447 = io_loadAddressDone_7 & _T_3446; // @[AxiStoreQueue.scala 143:36:@1634.4]
  assign noConflicts_7 = _T_3442 | _T_3447; // @[AxiStoreQueue.scala 142:95:@1635.4]
  assign _T_3450 = entriesToCheck_8 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1637.4]
  assign _T_3451 = _T_3450 | io_loadDataDone_8; // @[AxiStoreQueue.scala 142:64:@1638.4]
  assign _T_3455 = _GEN_911 != io_loadAddressQueue_8; // @[AxiStoreQueue.scala 143:56:@1639.4]
  assign _T_3456 = io_loadAddressDone_8 & _T_3455; // @[AxiStoreQueue.scala 143:36:@1640.4]
  assign noConflicts_8 = _T_3451 | _T_3456; // @[AxiStoreQueue.scala 142:95:@1641.4]
  assign _T_3459 = entriesToCheck_9 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1643.4]
  assign _T_3460 = _T_3459 | io_loadDataDone_9; // @[AxiStoreQueue.scala 142:64:@1644.4]
  assign _T_3464 = _GEN_911 != io_loadAddressQueue_9; // @[AxiStoreQueue.scala 143:56:@1645.4]
  assign _T_3465 = io_loadAddressDone_9 & _T_3464; // @[AxiStoreQueue.scala 143:36:@1646.4]
  assign noConflicts_9 = _T_3460 | _T_3465; // @[AxiStoreQueue.scala 142:95:@1647.4]
  assign _T_3468 = entriesToCheck_10 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1649.4]
  assign _T_3469 = _T_3468 | io_loadDataDone_10; // @[AxiStoreQueue.scala 142:64:@1650.4]
  assign _T_3473 = _GEN_911 != io_loadAddressQueue_10; // @[AxiStoreQueue.scala 143:56:@1651.4]
  assign _T_3474 = io_loadAddressDone_10 & _T_3473; // @[AxiStoreQueue.scala 143:36:@1652.4]
  assign noConflicts_10 = _T_3469 | _T_3474; // @[AxiStoreQueue.scala 142:95:@1653.4]
  assign _T_3477 = entriesToCheck_11 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1655.4]
  assign _T_3478 = _T_3477 | io_loadDataDone_11; // @[AxiStoreQueue.scala 142:64:@1656.4]
  assign _T_3482 = _GEN_911 != io_loadAddressQueue_11; // @[AxiStoreQueue.scala 143:56:@1657.4]
  assign _T_3483 = io_loadAddressDone_11 & _T_3482; // @[AxiStoreQueue.scala 143:36:@1658.4]
  assign noConflicts_11 = _T_3478 | _T_3483; // @[AxiStoreQueue.scala 142:95:@1659.4]
  assign _T_3486 = entriesToCheck_12 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1661.4]
  assign _T_3487 = _T_3486 | io_loadDataDone_12; // @[AxiStoreQueue.scala 142:64:@1662.4]
  assign _T_3491 = _GEN_911 != io_loadAddressQueue_12; // @[AxiStoreQueue.scala 143:56:@1663.4]
  assign _T_3492 = io_loadAddressDone_12 & _T_3491; // @[AxiStoreQueue.scala 143:36:@1664.4]
  assign noConflicts_12 = _T_3487 | _T_3492; // @[AxiStoreQueue.scala 142:95:@1665.4]
  assign _T_3495 = entriesToCheck_13 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1667.4]
  assign _T_3496 = _T_3495 | io_loadDataDone_13; // @[AxiStoreQueue.scala 142:64:@1668.4]
  assign _T_3500 = _GEN_911 != io_loadAddressQueue_13; // @[AxiStoreQueue.scala 143:56:@1669.4]
  assign _T_3501 = io_loadAddressDone_13 & _T_3500; // @[AxiStoreQueue.scala 143:36:@1670.4]
  assign noConflicts_13 = _T_3496 | _T_3501; // @[AxiStoreQueue.scala 142:95:@1671.4]
  assign _T_3504 = entriesToCheck_14 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1673.4]
  assign _T_3505 = _T_3504 | io_loadDataDone_14; // @[AxiStoreQueue.scala 142:64:@1674.4]
  assign _T_3509 = _GEN_911 != io_loadAddressQueue_14; // @[AxiStoreQueue.scala 143:56:@1675.4]
  assign _T_3510 = io_loadAddressDone_14 & _T_3509; // @[AxiStoreQueue.scala 143:36:@1676.4]
  assign noConflicts_14 = _T_3505 | _T_3510; // @[AxiStoreQueue.scala 142:95:@1677.4]
  assign _T_3513 = entriesToCheck_15 == 1'h0; // @[AxiStoreQueue.scala 142:34:@1679.4]
  assign _T_3514 = _T_3513 | io_loadDataDone_15; // @[AxiStoreQueue.scala 142:64:@1680.4]
  assign _T_3518 = _GEN_911 != io_loadAddressQueue_15; // @[AxiStoreQueue.scala 143:56:@1681.4]
  assign _T_3519 = io_loadAddressDone_15 & _T_3518; // @[AxiStoreQueue.scala 143:36:@1682.4]
  assign noConflicts_15 = _T_3514 | _T_3519; // @[AxiStoreQueue.scala 142:95:@1683.4]
  assign _GEN_913 = 4'h1 == dummyHead ? addrKnown_1 : addrKnown_0; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_914 = 4'h2 == dummyHead ? addrKnown_2 : _GEN_913; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_915 = 4'h3 == dummyHead ? addrKnown_3 : _GEN_914; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_916 = 4'h4 == dummyHead ? addrKnown_4 : _GEN_915; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_917 = 4'h5 == dummyHead ? addrKnown_5 : _GEN_916; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_918 = 4'h6 == dummyHead ? addrKnown_6 : _GEN_917; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_919 = 4'h7 == dummyHead ? addrKnown_7 : _GEN_918; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_920 = 4'h8 == dummyHead ? addrKnown_8 : _GEN_919; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_921 = 4'h9 == dummyHead ? addrKnown_9 : _GEN_920; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_922 = 4'ha == dummyHead ? addrKnown_10 : _GEN_921; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_923 = 4'hb == dummyHead ? addrKnown_11 : _GEN_922; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_924 = 4'hc == dummyHead ? addrKnown_12 : _GEN_923; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_925 = 4'hd == dummyHead ? addrKnown_13 : _GEN_924; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_926 = 4'he == dummyHead ? addrKnown_14 : _GEN_925; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_927 = 4'hf == dummyHead ? addrKnown_15 : _GEN_926; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_929 = 4'h1 == dummyHead ? dataKnown_1 : dataKnown_0; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_930 = 4'h2 == dummyHead ? dataKnown_2 : _GEN_929; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_931 = 4'h3 == dummyHead ? dataKnown_3 : _GEN_930; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_932 = 4'h4 == dummyHead ? dataKnown_4 : _GEN_931; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_933 = 4'h5 == dummyHead ? dataKnown_5 : _GEN_932; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_934 = 4'h6 == dummyHead ? dataKnown_6 : _GEN_933; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_935 = 4'h7 == dummyHead ? dataKnown_7 : _GEN_934; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_936 = 4'h8 == dummyHead ? dataKnown_8 : _GEN_935; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_937 = 4'h9 == dummyHead ? dataKnown_9 : _GEN_936; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_938 = 4'ha == dummyHead ? dataKnown_10 : _GEN_937; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_939 = 4'hb == dummyHead ? dataKnown_11 : _GEN_938; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_940 = 4'hc == dummyHead ? dataKnown_12 : _GEN_939; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_941 = 4'hd == dummyHead ? dataKnown_13 : _GEN_940; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_942 = 4'he == dummyHead ? dataKnown_14 : _GEN_941; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_943 = 4'hf == dummyHead ? dataKnown_15 : _GEN_942; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _T_3527 = _GEN_927 & _GEN_943; // @[AxiStoreQueue.scala 156:49:@1685.4]
  assign _GEN_945 = 4'h1 == dummyHead ? storeCompleted_1 : storeCompleted_0; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_946 = 4'h2 == dummyHead ? storeCompleted_2 : _GEN_945; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_947 = 4'h3 == dummyHead ? storeCompleted_3 : _GEN_946; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_948 = 4'h4 == dummyHead ? storeCompleted_4 : _GEN_947; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_949 = 4'h5 == dummyHead ? storeCompleted_5 : _GEN_948; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_950 = 4'h6 == dummyHead ? storeCompleted_6 : _GEN_949; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_951 = 4'h7 == dummyHead ? storeCompleted_7 : _GEN_950; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_952 = 4'h8 == dummyHead ? storeCompleted_8 : _GEN_951; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_953 = 4'h9 == dummyHead ? storeCompleted_9 : _GEN_952; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_954 = 4'ha == dummyHead ? storeCompleted_10 : _GEN_953; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_955 = 4'hb == dummyHead ? storeCompleted_11 : _GEN_954; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_956 = 4'hc == dummyHead ? storeCompleted_12 : _GEN_955; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_957 = 4'hd == dummyHead ? storeCompleted_13 : _GEN_956; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_958 = 4'he == dummyHead ? storeCompleted_14 : _GEN_957; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _GEN_959 = 4'hf == dummyHead ? storeCompleted_15 : _GEN_958; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _T_3532 = _GEN_959 == 1'h0; // @[AxiStoreQueue.scala 156:76:@1686.4]
  assign _T_3533 = _T_3527 & _T_3532; // @[AxiStoreQueue.scala 156:73:@1687.4]
  assign _T_3536 = noConflicts_0 & noConflicts_1; // @[AxiStoreQueue.scala 156:124:@1689.4]
  assign _T_3537 = _T_3536 & noConflicts_2; // @[AxiStoreQueue.scala 156:124:@1690.4]
  assign _T_3538 = _T_3537 & noConflicts_3; // @[AxiStoreQueue.scala 156:124:@1691.4]
  assign _T_3539 = _T_3538 & noConflicts_4; // @[AxiStoreQueue.scala 156:124:@1692.4]
  assign _T_3540 = _T_3539 & noConflicts_5; // @[AxiStoreQueue.scala 156:124:@1693.4]
  assign _T_3541 = _T_3540 & noConflicts_6; // @[AxiStoreQueue.scala 156:124:@1694.4]
  assign _T_3542 = _T_3541 & noConflicts_7; // @[AxiStoreQueue.scala 156:124:@1695.4]
  assign _T_3543 = _T_3542 & noConflicts_8; // @[AxiStoreQueue.scala 156:124:@1696.4]
  assign _T_3544 = _T_3543 & noConflicts_9; // @[AxiStoreQueue.scala 156:124:@1697.4]
  assign _T_3545 = _T_3544 & noConflicts_10; // @[AxiStoreQueue.scala 156:124:@1698.4]
  assign _T_3546 = _T_3545 & noConflicts_11; // @[AxiStoreQueue.scala 156:124:@1699.4]
  assign _T_3547 = _T_3546 & noConflicts_12; // @[AxiStoreQueue.scala 156:124:@1700.4]
  assign _T_3548 = _T_3547 & noConflicts_13; // @[AxiStoreQueue.scala 156:124:@1701.4]
  assign _T_3549 = _T_3548 & noConflicts_14; // @[AxiStoreQueue.scala 156:124:@1702.4]
  assign _T_3550 = _T_3549 & noConflicts_15; // @[AxiStoreQueue.scala 156:124:@1703.4]
  assign storeRequest = _T_3533 & _T_3550; // @[AxiStoreQueue.scala 156:103:@1704.4]
  assign _T_3553 = io_storeQIdxIn == 4'h0; // @[AxiStoreQueue.scala 168:54:@1710.6]
  assign _T_3554 = io_storeQIdxInValid & _T_3553; // @[AxiStoreQueue.scala 168:36:@1711.6]
  assign _GEN_960 = _T_3554 ? 1'h1 : storeCompleted_0; // @[AxiStoreQueue.scala 168:75:@1712.6]
  assign _GEN_961 = initBits_0 ? 1'h0 : _GEN_960; // @[AxiStoreQueue.scala 166:35:@1706.4]
  assign _T_3558 = io_storeQIdxIn == 4'h1; // @[AxiStoreQueue.scala 168:54:@1719.6]
  assign _T_3559 = io_storeQIdxInValid & _T_3558; // @[AxiStoreQueue.scala 168:36:@1720.6]
  assign _GEN_962 = _T_3559 ? 1'h1 : storeCompleted_1; // @[AxiStoreQueue.scala 168:75:@1721.6]
  assign _GEN_963 = initBits_1 ? 1'h0 : _GEN_962; // @[AxiStoreQueue.scala 166:35:@1715.4]
  assign _T_3563 = io_storeQIdxIn == 4'h2; // @[AxiStoreQueue.scala 168:54:@1728.6]
  assign _T_3564 = io_storeQIdxInValid & _T_3563; // @[AxiStoreQueue.scala 168:36:@1729.6]
  assign _GEN_964 = _T_3564 ? 1'h1 : storeCompleted_2; // @[AxiStoreQueue.scala 168:75:@1730.6]
  assign _GEN_965 = initBits_2 ? 1'h0 : _GEN_964; // @[AxiStoreQueue.scala 166:35:@1724.4]
  assign _T_3568 = io_storeQIdxIn == 4'h3; // @[AxiStoreQueue.scala 168:54:@1737.6]
  assign _T_3569 = io_storeQIdxInValid & _T_3568; // @[AxiStoreQueue.scala 168:36:@1738.6]
  assign _GEN_966 = _T_3569 ? 1'h1 : storeCompleted_3; // @[AxiStoreQueue.scala 168:75:@1739.6]
  assign _GEN_967 = initBits_3 ? 1'h0 : _GEN_966; // @[AxiStoreQueue.scala 166:35:@1733.4]
  assign _T_3573 = io_storeQIdxIn == 4'h4; // @[AxiStoreQueue.scala 168:54:@1746.6]
  assign _T_3574 = io_storeQIdxInValid & _T_3573; // @[AxiStoreQueue.scala 168:36:@1747.6]
  assign _GEN_968 = _T_3574 ? 1'h1 : storeCompleted_4; // @[AxiStoreQueue.scala 168:75:@1748.6]
  assign _GEN_969 = initBits_4 ? 1'h0 : _GEN_968; // @[AxiStoreQueue.scala 166:35:@1742.4]
  assign _T_3578 = io_storeQIdxIn == 4'h5; // @[AxiStoreQueue.scala 168:54:@1755.6]
  assign _T_3579 = io_storeQIdxInValid & _T_3578; // @[AxiStoreQueue.scala 168:36:@1756.6]
  assign _GEN_970 = _T_3579 ? 1'h1 : storeCompleted_5; // @[AxiStoreQueue.scala 168:75:@1757.6]
  assign _GEN_971 = initBits_5 ? 1'h0 : _GEN_970; // @[AxiStoreQueue.scala 166:35:@1751.4]
  assign _T_3583 = io_storeQIdxIn == 4'h6; // @[AxiStoreQueue.scala 168:54:@1764.6]
  assign _T_3584 = io_storeQIdxInValid & _T_3583; // @[AxiStoreQueue.scala 168:36:@1765.6]
  assign _GEN_972 = _T_3584 ? 1'h1 : storeCompleted_6; // @[AxiStoreQueue.scala 168:75:@1766.6]
  assign _GEN_973 = initBits_6 ? 1'h0 : _GEN_972; // @[AxiStoreQueue.scala 166:35:@1760.4]
  assign _T_3588 = io_storeQIdxIn == 4'h7; // @[AxiStoreQueue.scala 168:54:@1773.6]
  assign _T_3589 = io_storeQIdxInValid & _T_3588; // @[AxiStoreQueue.scala 168:36:@1774.6]
  assign _GEN_974 = _T_3589 ? 1'h1 : storeCompleted_7; // @[AxiStoreQueue.scala 168:75:@1775.6]
  assign _GEN_975 = initBits_7 ? 1'h0 : _GEN_974; // @[AxiStoreQueue.scala 166:35:@1769.4]
  assign _T_3593 = io_storeQIdxIn == 4'h8; // @[AxiStoreQueue.scala 168:54:@1782.6]
  assign _T_3594 = io_storeQIdxInValid & _T_3593; // @[AxiStoreQueue.scala 168:36:@1783.6]
  assign _GEN_976 = _T_3594 ? 1'h1 : storeCompleted_8; // @[AxiStoreQueue.scala 168:75:@1784.6]
  assign _GEN_977 = initBits_8 ? 1'h0 : _GEN_976; // @[AxiStoreQueue.scala 166:35:@1778.4]
  assign _T_3598 = io_storeQIdxIn == 4'h9; // @[AxiStoreQueue.scala 168:54:@1791.6]
  assign _T_3599 = io_storeQIdxInValid & _T_3598; // @[AxiStoreQueue.scala 168:36:@1792.6]
  assign _GEN_978 = _T_3599 ? 1'h1 : storeCompleted_9; // @[AxiStoreQueue.scala 168:75:@1793.6]
  assign _GEN_979 = initBits_9 ? 1'h0 : _GEN_978; // @[AxiStoreQueue.scala 166:35:@1787.4]
  assign _T_3603 = io_storeQIdxIn == 4'ha; // @[AxiStoreQueue.scala 168:54:@1800.6]
  assign _T_3604 = io_storeQIdxInValid & _T_3603; // @[AxiStoreQueue.scala 168:36:@1801.6]
  assign _GEN_980 = _T_3604 ? 1'h1 : storeCompleted_10; // @[AxiStoreQueue.scala 168:75:@1802.6]
  assign _GEN_981 = initBits_10 ? 1'h0 : _GEN_980; // @[AxiStoreQueue.scala 166:35:@1796.4]
  assign _T_3608 = io_storeQIdxIn == 4'hb; // @[AxiStoreQueue.scala 168:54:@1809.6]
  assign _T_3609 = io_storeQIdxInValid & _T_3608; // @[AxiStoreQueue.scala 168:36:@1810.6]
  assign _GEN_982 = _T_3609 ? 1'h1 : storeCompleted_11; // @[AxiStoreQueue.scala 168:75:@1811.6]
  assign _GEN_983 = initBits_11 ? 1'h0 : _GEN_982; // @[AxiStoreQueue.scala 166:35:@1805.4]
  assign _T_3613 = io_storeQIdxIn == 4'hc; // @[AxiStoreQueue.scala 168:54:@1818.6]
  assign _T_3614 = io_storeQIdxInValid & _T_3613; // @[AxiStoreQueue.scala 168:36:@1819.6]
  assign _GEN_984 = _T_3614 ? 1'h1 : storeCompleted_12; // @[AxiStoreQueue.scala 168:75:@1820.6]
  assign _GEN_985 = initBits_12 ? 1'h0 : _GEN_984; // @[AxiStoreQueue.scala 166:35:@1814.4]
  assign _T_3618 = io_storeQIdxIn == 4'hd; // @[AxiStoreQueue.scala 168:54:@1827.6]
  assign _T_3619 = io_storeQIdxInValid & _T_3618; // @[AxiStoreQueue.scala 168:36:@1828.6]
  assign _GEN_986 = _T_3619 ? 1'h1 : storeCompleted_13; // @[AxiStoreQueue.scala 168:75:@1829.6]
  assign _GEN_987 = initBits_13 ? 1'h0 : _GEN_986; // @[AxiStoreQueue.scala 166:35:@1823.4]
  assign _T_3623 = io_storeQIdxIn == 4'he; // @[AxiStoreQueue.scala 168:54:@1836.6]
  assign _T_3624 = io_storeQIdxInValid & _T_3623; // @[AxiStoreQueue.scala 168:36:@1837.6]
  assign _GEN_988 = _T_3624 ? 1'h1 : storeCompleted_14; // @[AxiStoreQueue.scala 168:75:@1838.6]
  assign _GEN_989 = initBits_14 ? 1'h0 : _GEN_988; // @[AxiStoreQueue.scala 166:35:@1832.4]
  assign _T_3628 = io_storeQIdxIn == 4'hf; // @[AxiStoreQueue.scala 168:54:@1845.6]
  assign _T_3629 = io_storeQIdxInValid & _T_3628; // @[AxiStoreQueue.scala 168:36:@1846.6]
  assign _GEN_990 = _T_3629 ? 1'h1 : storeCompleted_15; // @[AxiStoreQueue.scala 168:75:@1847.6]
  assign _GEN_991 = initBits_15 ? 1'h0 : _GEN_990; // @[AxiStoreQueue.scala 166:35:@1841.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1851.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1853.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1855.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1857.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1859.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1861.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1863.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1865.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1867.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1869.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1871.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1873.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1875.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1877.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1879.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[AxiStoreQueue.scala 185:72:@1881.4]
  assign _T_4114 = addrKnown_0 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1885.4]
  assign _T_4115 = entriesPorts_0_0 & _T_4114; // @[AxiStoreQueue.scala 197:88:@1886.4]
  assign _T_4117 = addrKnown_1 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1887.4]
  assign _T_4118 = entriesPorts_0_1 & _T_4117; // @[AxiStoreQueue.scala 197:88:@1888.4]
  assign _T_4120 = addrKnown_2 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1889.4]
  assign _T_4121 = entriesPorts_0_2 & _T_4120; // @[AxiStoreQueue.scala 197:88:@1890.4]
  assign _T_4123 = addrKnown_3 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1891.4]
  assign _T_4124 = entriesPorts_0_3 & _T_4123; // @[AxiStoreQueue.scala 197:88:@1892.4]
  assign _T_4126 = addrKnown_4 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1893.4]
  assign _T_4127 = entriesPorts_0_4 & _T_4126; // @[AxiStoreQueue.scala 197:88:@1894.4]
  assign _T_4129 = addrKnown_5 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1895.4]
  assign _T_4130 = entriesPorts_0_5 & _T_4129; // @[AxiStoreQueue.scala 197:88:@1896.4]
  assign _T_4132 = addrKnown_6 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1897.4]
  assign _T_4133 = entriesPorts_0_6 & _T_4132; // @[AxiStoreQueue.scala 197:88:@1898.4]
  assign _T_4135 = addrKnown_7 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1899.4]
  assign _T_4136 = entriesPorts_0_7 & _T_4135; // @[AxiStoreQueue.scala 197:88:@1900.4]
  assign _T_4138 = addrKnown_8 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1901.4]
  assign _T_4139 = entriesPorts_0_8 & _T_4138; // @[AxiStoreQueue.scala 197:88:@1902.4]
  assign _T_4141 = addrKnown_9 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1903.4]
  assign _T_4142 = entriesPorts_0_9 & _T_4141; // @[AxiStoreQueue.scala 197:88:@1904.4]
  assign _T_4144 = addrKnown_10 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1905.4]
  assign _T_4145 = entriesPorts_0_10 & _T_4144; // @[AxiStoreQueue.scala 197:88:@1906.4]
  assign _T_4147 = addrKnown_11 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1907.4]
  assign _T_4148 = entriesPorts_0_11 & _T_4147; // @[AxiStoreQueue.scala 197:88:@1908.4]
  assign _T_4150 = addrKnown_12 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1909.4]
  assign _T_4151 = entriesPorts_0_12 & _T_4150; // @[AxiStoreQueue.scala 197:88:@1910.4]
  assign _T_4153 = addrKnown_13 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1911.4]
  assign _T_4154 = entriesPorts_0_13 & _T_4153; // @[AxiStoreQueue.scala 197:88:@1912.4]
  assign _T_4156 = addrKnown_14 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1913.4]
  assign _T_4157 = entriesPorts_0_14 & _T_4156; // @[AxiStoreQueue.scala 197:88:@1914.4]
  assign _T_4159 = addrKnown_15 == 1'h0; // @[AxiStoreQueue.scala 197:91:@1915.4]
  assign _T_4160 = entriesPorts_0_15 & _T_4159; // @[AxiStoreQueue.scala 197:88:@1916.4]
  assign _T_4184 = dataKnown_0 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1934.4]
  assign _T_4185 = entriesPorts_0_0 & _T_4184; // @[AxiStoreQueue.scala 198:88:@1935.4]
  assign _T_4187 = dataKnown_1 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1936.4]
  assign _T_4188 = entriesPorts_0_1 & _T_4187; // @[AxiStoreQueue.scala 198:88:@1937.4]
  assign _T_4190 = dataKnown_2 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1938.4]
  assign _T_4191 = entriesPorts_0_2 & _T_4190; // @[AxiStoreQueue.scala 198:88:@1939.4]
  assign _T_4193 = dataKnown_3 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1940.4]
  assign _T_4194 = entriesPorts_0_3 & _T_4193; // @[AxiStoreQueue.scala 198:88:@1941.4]
  assign _T_4196 = dataKnown_4 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1942.4]
  assign _T_4197 = entriesPorts_0_4 & _T_4196; // @[AxiStoreQueue.scala 198:88:@1943.4]
  assign _T_4199 = dataKnown_5 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1944.4]
  assign _T_4200 = entriesPorts_0_5 & _T_4199; // @[AxiStoreQueue.scala 198:88:@1945.4]
  assign _T_4202 = dataKnown_6 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1946.4]
  assign _T_4203 = entriesPorts_0_6 & _T_4202; // @[AxiStoreQueue.scala 198:88:@1947.4]
  assign _T_4205 = dataKnown_7 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1948.4]
  assign _T_4206 = entriesPorts_0_7 & _T_4205; // @[AxiStoreQueue.scala 198:88:@1949.4]
  assign _T_4208 = dataKnown_8 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1950.4]
  assign _T_4209 = entriesPorts_0_8 & _T_4208; // @[AxiStoreQueue.scala 198:88:@1951.4]
  assign _T_4211 = dataKnown_9 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1952.4]
  assign _T_4212 = entriesPorts_0_9 & _T_4211; // @[AxiStoreQueue.scala 198:88:@1953.4]
  assign _T_4214 = dataKnown_10 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1954.4]
  assign _T_4215 = entriesPorts_0_10 & _T_4214; // @[AxiStoreQueue.scala 198:88:@1955.4]
  assign _T_4217 = dataKnown_11 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1956.4]
  assign _T_4218 = entriesPorts_0_11 & _T_4217; // @[AxiStoreQueue.scala 198:88:@1957.4]
  assign _T_4220 = dataKnown_12 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1958.4]
  assign _T_4221 = entriesPorts_0_12 & _T_4220; // @[AxiStoreQueue.scala 198:88:@1959.4]
  assign _T_4223 = dataKnown_13 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1960.4]
  assign _T_4224 = entriesPorts_0_13 & _T_4223; // @[AxiStoreQueue.scala 198:88:@1961.4]
  assign _T_4226 = dataKnown_14 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1962.4]
  assign _T_4227 = entriesPorts_0_14 & _T_4226; // @[AxiStoreQueue.scala 198:88:@1963.4]
  assign _T_4229 = dataKnown_15 == 1'h0; // @[AxiStoreQueue.scala 198:91:@1964.4]
  assign _T_4230 = entriesPorts_0_15 & _T_4229; // @[AxiStoreQueue.scala 198:88:@1965.4]
  assign _T_4255 = 16'h1 << dummyHead; // @[OneHot.scala 52:12:@1984.4]
  assign _T_4257 = _T_4255[0]; // @[util.scala 33:60:@1986.4]
  assign _T_4258 = _T_4255[1]; // @[util.scala 33:60:@1987.4]
  assign _T_4259 = _T_4255[2]; // @[util.scala 33:60:@1988.4]
  assign _T_4260 = _T_4255[3]; // @[util.scala 33:60:@1989.4]
  assign _T_4261 = _T_4255[4]; // @[util.scala 33:60:@1990.4]
  assign _T_4262 = _T_4255[5]; // @[util.scala 33:60:@1991.4]
  assign _T_4263 = _T_4255[6]; // @[util.scala 33:60:@1992.4]
  assign _T_4264 = _T_4255[7]; // @[util.scala 33:60:@1993.4]
  assign _T_4265 = _T_4255[8]; // @[util.scala 33:60:@1994.4]
  assign _T_4266 = _T_4255[9]; // @[util.scala 33:60:@1995.4]
  assign _T_4267 = _T_4255[10]; // @[util.scala 33:60:@1996.4]
  assign _T_4268 = _T_4255[11]; // @[util.scala 33:60:@1997.4]
  assign _T_4269 = _T_4255[12]; // @[util.scala 33:60:@1998.4]
  assign _T_4270 = _T_4255[13]; // @[util.scala 33:60:@1999.4]
  assign _T_4271 = _T_4255[14]; // @[util.scala 33:60:@2000.4]
  assign _T_4272 = _T_4255[15]; // @[util.scala 33:60:@2001.4]
  assign _T_4313 = _T_4160 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2019.4]
  assign _T_4314 = _T_4157 ? 16'h4000 : _T_4313; // @[Mux.scala 31:69:@2020.4]
  assign _T_4315 = _T_4154 ? 16'h2000 : _T_4314; // @[Mux.scala 31:69:@2021.4]
  assign _T_4316 = _T_4151 ? 16'h1000 : _T_4315; // @[Mux.scala 31:69:@2022.4]
  assign _T_4317 = _T_4148 ? 16'h800 : _T_4316; // @[Mux.scala 31:69:@2023.4]
  assign _T_4318 = _T_4145 ? 16'h400 : _T_4317; // @[Mux.scala 31:69:@2024.4]
  assign _T_4319 = _T_4142 ? 16'h200 : _T_4318; // @[Mux.scala 31:69:@2025.4]
  assign _T_4320 = _T_4139 ? 16'h100 : _T_4319; // @[Mux.scala 31:69:@2026.4]
  assign _T_4321 = _T_4136 ? 16'h80 : _T_4320; // @[Mux.scala 31:69:@2027.4]
  assign _T_4322 = _T_4133 ? 16'h40 : _T_4321; // @[Mux.scala 31:69:@2028.4]
  assign _T_4323 = _T_4130 ? 16'h20 : _T_4322; // @[Mux.scala 31:69:@2029.4]
  assign _T_4324 = _T_4127 ? 16'h10 : _T_4323; // @[Mux.scala 31:69:@2030.4]
  assign _T_4325 = _T_4124 ? 16'h8 : _T_4324; // @[Mux.scala 31:69:@2031.4]
  assign _T_4326 = _T_4121 ? 16'h4 : _T_4325; // @[Mux.scala 31:69:@2032.4]
  assign _T_4327 = _T_4118 ? 16'h2 : _T_4326; // @[Mux.scala 31:69:@2033.4]
  assign _T_4328 = _T_4115 ? 16'h1 : _T_4327; // @[Mux.scala 31:69:@2034.4]
  assign _T_4329 = _T_4328[0]; // @[OneHot.scala 66:30:@2035.4]
  assign _T_4330 = _T_4328[1]; // @[OneHot.scala 66:30:@2036.4]
  assign _T_4331 = _T_4328[2]; // @[OneHot.scala 66:30:@2037.4]
  assign _T_4332 = _T_4328[3]; // @[OneHot.scala 66:30:@2038.4]
  assign _T_4333 = _T_4328[4]; // @[OneHot.scala 66:30:@2039.4]
  assign _T_4334 = _T_4328[5]; // @[OneHot.scala 66:30:@2040.4]
  assign _T_4335 = _T_4328[6]; // @[OneHot.scala 66:30:@2041.4]
  assign _T_4336 = _T_4328[7]; // @[OneHot.scala 66:30:@2042.4]
  assign _T_4337 = _T_4328[8]; // @[OneHot.scala 66:30:@2043.4]
  assign _T_4338 = _T_4328[9]; // @[OneHot.scala 66:30:@2044.4]
  assign _T_4339 = _T_4328[10]; // @[OneHot.scala 66:30:@2045.4]
  assign _T_4340 = _T_4328[11]; // @[OneHot.scala 66:30:@2046.4]
  assign _T_4341 = _T_4328[12]; // @[OneHot.scala 66:30:@2047.4]
  assign _T_4342 = _T_4328[13]; // @[OneHot.scala 66:30:@2048.4]
  assign _T_4343 = _T_4328[14]; // @[OneHot.scala 66:30:@2049.4]
  assign _T_4344 = _T_4328[15]; // @[OneHot.scala 66:30:@2050.4]
  assign _T_4385 = _T_4115 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2068.4]
  assign _T_4386 = _T_4160 ? 16'h4000 : _T_4385; // @[Mux.scala 31:69:@2069.4]
  assign _T_4387 = _T_4157 ? 16'h2000 : _T_4386; // @[Mux.scala 31:69:@2070.4]
  assign _T_4388 = _T_4154 ? 16'h1000 : _T_4387; // @[Mux.scala 31:69:@2071.4]
  assign _T_4389 = _T_4151 ? 16'h800 : _T_4388; // @[Mux.scala 31:69:@2072.4]
  assign _T_4390 = _T_4148 ? 16'h400 : _T_4389; // @[Mux.scala 31:69:@2073.4]
  assign _T_4391 = _T_4145 ? 16'h200 : _T_4390; // @[Mux.scala 31:69:@2074.4]
  assign _T_4392 = _T_4142 ? 16'h100 : _T_4391; // @[Mux.scala 31:69:@2075.4]
  assign _T_4393 = _T_4139 ? 16'h80 : _T_4392; // @[Mux.scala 31:69:@2076.4]
  assign _T_4394 = _T_4136 ? 16'h40 : _T_4393; // @[Mux.scala 31:69:@2077.4]
  assign _T_4395 = _T_4133 ? 16'h20 : _T_4394; // @[Mux.scala 31:69:@2078.4]
  assign _T_4396 = _T_4130 ? 16'h10 : _T_4395; // @[Mux.scala 31:69:@2079.4]
  assign _T_4397 = _T_4127 ? 16'h8 : _T_4396; // @[Mux.scala 31:69:@2080.4]
  assign _T_4398 = _T_4124 ? 16'h4 : _T_4397; // @[Mux.scala 31:69:@2081.4]
  assign _T_4399 = _T_4121 ? 16'h2 : _T_4398; // @[Mux.scala 31:69:@2082.4]
  assign _T_4400 = _T_4118 ? 16'h1 : _T_4399; // @[Mux.scala 31:69:@2083.4]
  assign _T_4401 = _T_4400[0]; // @[OneHot.scala 66:30:@2084.4]
  assign _T_4402 = _T_4400[1]; // @[OneHot.scala 66:30:@2085.4]
  assign _T_4403 = _T_4400[2]; // @[OneHot.scala 66:30:@2086.4]
  assign _T_4404 = _T_4400[3]; // @[OneHot.scala 66:30:@2087.4]
  assign _T_4405 = _T_4400[4]; // @[OneHot.scala 66:30:@2088.4]
  assign _T_4406 = _T_4400[5]; // @[OneHot.scala 66:30:@2089.4]
  assign _T_4407 = _T_4400[6]; // @[OneHot.scala 66:30:@2090.4]
  assign _T_4408 = _T_4400[7]; // @[OneHot.scala 66:30:@2091.4]
  assign _T_4409 = _T_4400[8]; // @[OneHot.scala 66:30:@2092.4]
  assign _T_4410 = _T_4400[9]; // @[OneHot.scala 66:30:@2093.4]
  assign _T_4411 = _T_4400[10]; // @[OneHot.scala 66:30:@2094.4]
  assign _T_4412 = _T_4400[11]; // @[OneHot.scala 66:30:@2095.4]
  assign _T_4413 = _T_4400[12]; // @[OneHot.scala 66:30:@2096.4]
  assign _T_4414 = _T_4400[13]; // @[OneHot.scala 66:30:@2097.4]
  assign _T_4415 = _T_4400[14]; // @[OneHot.scala 66:30:@2098.4]
  assign _T_4416 = _T_4400[15]; // @[OneHot.scala 66:30:@2099.4]
  assign _T_4457 = _T_4118 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2117.4]
  assign _T_4458 = _T_4115 ? 16'h4000 : _T_4457; // @[Mux.scala 31:69:@2118.4]
  assign _T_4459 = _T_4160 ? 16'h2000 : _T_4458; // @[Mux.scala 31:69:@2119.4]
  assign _T_4460 = _T_4157 ? 16'h1000 : _T_4459; // @[Mux.scala 31:69:@2120.4]
  assign _T_4461 = _T_4154 ? 16'h800 : _T_4460; // @[Mux.scala 31:69:@2121.4]
  assign _T_4462 = _T_4151 ? 16'h400 : _T_4461; // @[Mux.scala 31:69:@2122.4]
  assign _T_4463 = _T_4148 ? 16'h200 : _T_4462; // @[Mux.scala 31:69:@2123.4]
  assign _T_4464 = _T_4145 ? 16'h100 : _T_4463; // @[Mux.scala 31:69:@2124.4]
  assign _T_4465 = _T_4142 ? 16'h80 : _T_4464; // @[Mux.scala 31:69:@2125.4]
  assign _T_4466 = _T_4139 ? 16'h40 : _T_4465; // @[Mux.scala 31:69:@2126.4]
  assign _T_4467 = _T_4136 ? 16'h20 : _T_4466; // @[Mux.scala 31:69:@2127.4]
  assign _T_4468 = _T_4133 ? 16'h10 : _T_4467; // @[Mux.scala 31:69:@2128.4]
  assign _T_4469 = _T_4130 ? 16'h8 : _T_4468; // @[Mux.scala 31:69:@2129.4]
  assign _T_4470 = _T_4127 ? 16'h4 : _T_4469; // @[Mux.scala 31:69:@2130.4]
  assign _T_4471 = _T_4124 ? 16'h2 : _T_4470; // @[Mux.scala 31:69:@2131.4]
  assign _T_4472 = _T_4121 ? 16'h1 : _T_4471; // @[Mux.scala 31:69:@2132.4]
  assign _T_4473 = _T_4472[0]; // @[OneHot.scala 66:30:@2133.4]
  assign _T_4474 = _T_4472[1]; // @[OneHot.scala 66:30:@2134.4]
  assign _T_4475 = _T_4472[2]; // @[OneHot.scala 66:30:@2135.4]
  assign _T_4476 = _T_4472[3]; // @[OneHot.scala 66:30:@2136.4]
  assign _T_4477 = _T_4472[4]; // @[OneHot.scala 66:30:@2137.4]
  assign _T_4478 = _T_4472[5]; // @[OneHot.scala 66:30:@2138.4]
  assign _T_4479 = _T_4472[6]; // @[OneHot.scala 66:30:@2139.4]
  assign _T_4480 = _T_4472[7]; // @[OneHot.scala 66:30:@2140.4]
  assign _T_4481 = _T_4472[8]; // @[OneHot.scala 66:30:@2141.4]
  assign _T_4482 = _T_4472[9]; // @[OneHot.scala 66:30:@2142.4]
  assign _T_4483 = _T_4472[10]; // @[OneHot.scala 66:30:@2143.4]
  assign _T_4484 = _T_4472[11]; // @[OneHot.scala 66:30:@2144.4]
  assign _T_4485 = _T_4472[12]; // @[OneHot.scala 66:30:@2145.4]
  assign _T_4486 = _T_4472[13]; // @[OneHot.scala 66:30:@2146.4]
  assign _T_4487 = _T_4472[14]; // @[OneHot.scala 66:30:@2147.4]
  assign _T_4488 = _T_4472[15]; // @[OneHot.scala 66:30:@2148.4]
  assign _T_4529 = _T_4121 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2166.4]
  assign _T_4530 = _T_4118 ? 16'h4000 : _T_4529; // @[Mux.scala 31:69:@2167.4]
  assign _T_4531 = _T_4115 ? 16'h2000 : _T_4530; // @[Mux.scala 31:69:@2168.4]
  assign _T_4532 = _T_4160 ? 16'h1000 : _T_4531; // @[Mux.scala 31:69:@2169.4]
  assign _T_4533 = _T_4157 ? 16'h800 : _T_4532; // @[Mux.scala 31:69:@2170.4]
  assign _T_4534 = _T_4154 ? 16'h400 : _T_4533; // @[Mux.scala 31:69:@2171.4]
  assign _T_4535 = _T_4151 ? 16'h200 : _T_4534; // @[Mux.scala 31:69:@2172.4]
  assign _T_4536 = _T_4148 ? 16'h100 : _T_4535; // @[Mux.scala 31:69:@2173.4]
  assign _T_4537 = _T_4145 ? 16'h80 : _T_4536; // @[Mux.scala 31:69:@2174.4]
  assign _T_4538 = _T_4142 ? 16'h40 : _T_4537; // @[Mux.scala 31:69:@2175.4]
  assign _T_4539 = _T_4139 ? 16'h20 : _T_4538; // @[Mux.scala 31:69:@2176.4]
  assign _T_4540 = _T_4136 ? 16'h10 : _T_4539; // @[Mux.scala 31:69:@2177.4]
  assign _T_4541 = _T_4133 ? 16'h8 : _T_4540; // @[Mux.scala 31:69:@2178.4]
  assign _T_4542 = _T_4130 ? 16'h4 : _T_4541; // @[Mux.scala 31:69:@2179.4]
  assign _T_4543 = _T_4127 ? 16'h2 : _T_4542; // @[Mux.scala 31:69:@2180.4]
  assign _T_4544 = _T_4124 ? 16'h1 : _T_4543; // @[Mux.scala 31:69:@2181.4]
  assign _T_4545 = _T_4544[0]; // @[OneHot.scala 66:30:@2182.4]
  assign _T_4546 = _T_4544[1]; // @[OneHot.scala 66:30:@2183.4]
  assign _T_4547 = _T_4544[2]; // @[OneHot.scala 66:30:@2184.4]
  assign _T_4548 = _T_4544[3]; // @[OneHot.scala 66:30:@2185.4]
  assign _T_4549 = _T_4544[4]; // @[OneHot.scala 66:30:@2186.4]
  assign _T_4550 = _T_4544[5]; // @[OneHot.scala 66:30:@2187.4]
  assign _T_4551 = _T_4544[6]; // @[OneHot.scala 66:30:@2188.4]
  assign _T_4552 = _T_4544[7]; // @[OneHot.scala 66:30:@2189.4]
  assign _T_4553 = _T_4544[8]; // @[OneHot.scala 66:30:@2190.4]
  assign _T_4554 = _T_4544[9]; // @[OneHot.scala 66:30:@2191.4]
  assign _T_4555 = _T_4544[10]; // @[OneHot.scala 66:30:@2192.4]
  assign _T_4556 = _T_4544[11]; // @[OneHot.scala 66:30:@2193.4]
  assign _T_4557 = _T_4544[12]; // @[OneHot.scala 66:30:@2194.4]
  assign _T_4558 = _T_4544[13]; // @[OneHot.scala 66:30:@2195.4]
  assign _T_4559 = _T_4544[14]; // @[OneHot.scala 66:30:@2196.4]
  assign _T_4560 = _T_4544[15]; // @[OneHot.scala 66:30:@2197.4]
  assign _T_4601 = _T_4124 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2215.4]
  assign _T_4602 = _T_4121 ? 16'h4000 : _T_4601; // @[Mux.scala 31:69:@2216.4]
  assign _T_4603 = _T_4118 ? 16'h2000 : _T_4602; // @[Mux.scala 31:69:@2217.4]
  assign _T_4604 = _T_4115 ? 16'h1000 : _T_4603; // @[Mux.scala 31:69:@2218.4]
  assign _T_4605 = _T_4160 ? 16'h800 : _T_4604; // @[Mux.scala 31:69:@2219.4]
  assign _T_4606 = _T_4157 ? 16'h400 : _T_4605; // @[Mux.scala 31:69:@2220.4]
  assign _T_4607 = _T_4154 ? 16'h200 : _T_4606; // @[Mux.scala 31:69:@2221.4]
  assign _T_4608 = _T_4151 ? 16'h100 : _T_4607; // @[Mux.scala 31:69:@2222.4]
  assign _T_4609 = _T_4148 ? 16'h80 : _T_4608; // @[Mux.scala 31:69:@2223.4]
  assign _T_4610 = _T_4145 ? 16'h40 : _T_4609; // @[Mux.scala 31:69:@2224.4]
  assign _T_4611 = _T_4142 ? 16'h20 : _T_4610; // @[Mux.scala 31:69:@2225.4]
  assign _T_4612 = _T_4139 ? 16'h10 : _T_4611; // @[Mux.scala 31:69:@2226.4]
  assign _T_4613 = _T_4136 ? 16'h8 : _T_4612; // @[Mux.scala 31:69:@2227.4]
  assign _T_4614 = _T_4133 ? 16'h4 : _T_4613; // @[Mux.scala 31:69:@2228.4]
  assign _T_4615 = _T_4130 ? 16'h2 : _T_4614; // @[Mux.scala 31:69:@2229.4]
  assign _T_4616 = _T_4127 ? 16'h1 : _T_4615; // @[Mux.scala 31:69:@2230.4]
  assign _T_4617 = _T_4616[0]; // @[OneHot.scala 66:30:@2231.4]
  assign _T_4618 = _T_4616[1]; // @[OneHot.scala 66:30:@2232.4]
  assign _T_4619 = _T_4616[2]; // @[OneHot.scala 66:30:@2233.4]
  assign _T_4620 = _T_4616[3]; // @[OneHot.scala 66:30:@2234.4]
  assign _T_4621 = _T_4616[4]; // @[OneHot.scala 66:30:@2235.4]
  assign _T_4622 = _T_4616[5]; // @[OneHot.scala 66:30:@2236.4]
  assign _T_4623 = _T_4616[6]; // @[OneHot.scala 66:30:@2237.4]
  assign _T_4624 = _T_4616[7]; // @[OneHot.scala 66:30:@2238.4]
  assign _T_4625 = _T_4616[8]; // @[OneHot.scala 66:30:@2239.4]
  assign _T_4626 = _T_4616[9]; // @[OneHot.scala 66:30:@2240.4]
  assign _T_4627 = _T_4616[10]; // @[OneHot.scala 66:30:@2241.4]
  assign _T_4628 = _T_4616[11]; // @[OneHot.scala 66:30:@2242.4]
  assign _T_4629 = _T_4616[12]; // @[OneHot.scala 66:30:@2243.4]
  assign _T_4630 = _T_4616[13]; // @[OneHot.scala 66:30:@2244.4]
  assign _T_4631 = _T_4616[14]; // @[OneHot.scala 66:30:@2245.4]
  assign _T_4632 = _T_4616[15]; // @[OneHot.scala 66:30:@2246.4]
  assign _T_4673 = _T_4127 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2264.4]
  assign _T_4674 = _T_4124 ? 16'h4000 : _T_4673; // @[Mux.scala 31:69:@2265.4]
  assign _T_4675 = _T_4121 ? 16'h2000 : _T_4674; // @[Mux.scala 31:69:@2266.4]
  assign _T_4676 = _T_4118 ? 16'h1000 : _T_4675; // @[Mux.scala 31:69:@2267.4]
  assign _T_4677 = _T_4115 ? 16'h800 : _T_4676; // @[Mux.scala 31:69:@2268.4]
  assign _T_4678 = _T_4160 ? 16'h400 : _T_4677; // @[Mux.scala 31:69:@2269.4]
  assign _T_4679 = _T_4157 ? 16'h200 : _T_4678; // @[Mux.scala 31:69:@2270.4]
  assign _T_4680 = _T_4154 ? 16'h100 : _T_4679; // @[Mux.scala 31:69:@2271.4]
  assign _T_4681 = _T_4151 ? 16'h80 : _T_4680; // @[Mux.scala 31:69:@2272.4]
  assign _T_4682 = _T_4148 ? 16'h40 : _T_4681; // @[Mux.scala 31:69:@2273.4]
  assign _T_4683 = _T_4145 ? 16'h20 : _T_4682; // @[Mux.scala 31:69:@2274.4]
  assign _T_4684 = _T_4142 ? 16'h10 : _T_4683; // @[Mux.scala 31:69:@2275.4]
  assign _T_4685 = _T_4139 ? 16'h8 : _T_4684; // @[Mux.scala 31:69:@2276.4]
  assign _T_4686 = _T_4136 ? 16'h4 : _T_4685; // @[Mux.scala 31:69:@2277.4]
  assign _T_4687 = _T_4133 ? 16'h2 : _T_4686; // @[Mux.scala 31:69:@2278.4]
  assign _T_4688 = _T_4130 ? 16'h1 : _T_4687; // @[Mux.scala 31:69:@2279.4]
  assign _T_4689 = _T_4688[0]; // @[OneHot.scala 66:30:@2280.4]
  assign _T_4690 = _T_4688[1]; // @[OneHot.scala 66:30:@2281.4]
  assign _T_4691 = _T_4688[2]; // @[OneHot.scala 66:30:@2282.4]
  assign _T_4692 = _T_4688[3]; // @[OneHot.scala 66:30:@2283.4]
  assign _T_4693 = _T_4688[4]; // @[OneHot.scala 66:30:@2284.4]
  assign _T_4694 = _T_4688[5]; // @[OneHot.scala 66:30:@2285.4]
  assign _T_4695 = _T_4688[6]; // @[OneHot.scala 66:30:@2286.4]
  assign _T_4696 = _T_4688[7]; // @[OneHot.scala 66:30:@2287.4]
  assign _T_4697 = _T_4688[8]; // @[OneHot.scala 66:30:@2288.4]
  assign _T_4698 = _T_4688[9]; // @[OneHot.scala 66:30:@2289.4]
  assign _T_4699 = _T_4688[10]; // @[OneHot.scala 66:30:@2290.4]
  assign _T_4700 = _T_4688[11]; // @[OneHot.scala 66:30:@2291.4]
  assign _T_4701 = _T_4688[12]; // @[OneHot.scala 66:30:@2292.4]
  assign _T_4702 = _T_4688[13]; // @[OneHot.scala 66:30:@2293.4]
  assign _T_4703 = _T_4688[14]; // @[OneHot.scala 66:30:@2294.4]
  assign _T_4704 = _T_4688[15]; // @[OneHot.scala 66:30:@2295.4]
  assign _T_4745 = _T_4130 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2313.4]
  assign _T_4746 = _T_4127 ? 16'h4000 : _T_4745; // @[Mux.scala 31:69:@2314.4]
  assign _T_4747 = _T_4124 ? 16'h2000 : _T_4746; // @[Mux.scala 31:69:@2315.4]
  assign _T_4748 = _T_4121 ? 16'h1000 : _T_4747; // @[Mux.scala 31:69:@2316.4]
  assign _T_4749 = _T_4118 ? 16'h800 : _T_4748; // @[Mux.scala 31:69:@2317.4]
  assign _T_4750 = _T_4115 ? 16'h400 : _T_4749; // @[Mux.scala 31:69:@2318.4]
  assign _T_4751 = _T_4160 ? 16'h200 : _T_4750; // @[Mux.scala 31:69:@2319.4]
  assign _T_4752 = _T_4157 ? 16'h100 : _T_4751; // @[Mux.scala 31:69:@2320.4]
  assign _T_4753 = _T_4154 ? 16'h80 : _T_4752; // @[Mux.scala 31:69:@2321.4]
  assign _T_4754 = _T_4151 ? 16'h40 : _T_4753; // @[Mux.scala 31:69:@2322.4]
  assign _T_4755 = _T_4148 ? 16'h20 : _T_4754; // @[Mux.scala 31:69:@2323.4]
  assign _T_4756 = _T_4145 ? 16'h10 : _T_4755; // @[Mux.scala 31:69:@2324.4]
  assign _T_4757 = _T_4142 ? 16'h8 : _T_4756; // @[Mux.scala 31:69:@2325.4]
  assign _T_4758 = _T_4139 ? 16'h4 : _T_4757; // @[Mux.scala 31:69:@2326.4]
  assign _T_4759 = _T_4136 ? 16'h2 : _T_4758; // @[Mux.scala 31:69:@2327.4]
  assign _T_4760 = _T_4133 ? 16'h1 : _T_4759; // @[Mux.scala 31:69:@2328.4]
  assign _T_4761 = _T_4760[0]; // @[OneHot.scala 66:30:@2329.4]
  assign _T_4762 = _T_4760[1]; // @[OneHot.scala 66:30:@2330.4]
  assign _T_4763 = _T_4760[2]; // @[OneHot.scala 66:30:@2331.4]
  assign _T_4764 = _T_4760[3]; // @[OneHot.scala 66:30:@2332.4]
  assign _T_4765 = _T_4760[4]; // @[OneHot.scala 66:30:@2333.4]
  assign _T_4766 = _T_4760[5]; // @[OneHot.scala 66:30:@2334.4]
  assign _T_4767 = _T_4760[6]; // @[OneHot.scala 66:30:@2335.4]
  assign _T_4768 = _T_4760[7]; // @[OneHot.scala 66:30:@2336.4]
  assign _T_4769 = _T_4760[8]; // @[OneHot.scala 66:30:@2337.4]
  assign _T_4770 = _T_4760[9]; // @[OneHot.scala 66:30:@2338.4]
  assign _T_4771 = _T_4760[10]; // @[OneHot.scala 66:30:@2339.4]
  assign _T_4772 = _T_4760[11]; // @[OneHot.scala 66:30:@2340.4]
  assign _T_4773 = _T_4760[12]; // @[OneHot.scala 66:30:@2341.4]
  assign _T_4774 = _T_4760[13]; // @[OneHot.scala 66:30:@2342.4]
  assign _T_4775 = _T_4760[14]; // @[OneHot.scala 66:30:@2343.4]
  assign _T_4776 = _T_4760[15]; // @[OneHot.scala 66:30:@2344.4]
  assign _T_4817 = _T_4133 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2362.4]
  assign _T_4818 = _T_4130 ? 16'h4000 : _T_4817; // @[Mux.scala 31:69:@2363.4]
  assign _T_4819 = _T_4127 ? 16'h2000 : _T_4818; // @[Mux.scala 31:69:@2364.4]
  assign _T_4820 = _T_4124 ? 16'h1000 : _T_4819; // @[Mux.scala 31:69:@2365.4]
  assign _T_4821 = _T_4121 ? 16'h800 : _T_4820; // @[Mux.scala 31:69:@2366.4]
  assign _T_4822 = _T_4118 ? 16'h400 : _T_4821; // @[Mux.scala 31:69:@2367.4]
  assign _T_4823 = _T_4115 ? 16'h200 : _T_4822; // @[Mux.scala 31:69:@2368.4]
  assign _T_4824 = _T_4160 ? 16'h100 : _T_4823; // @[Mux.scala 31:69:@2369.4]
  assign _T_4825 = _T_4157 ? 16'h80 : _T_4824; // @[Mux.scala 31:69:@2370.4]
  assign _T_4826 = _T_4154 ? 16'h40 : _T_4825; // @[Mux.scala 31:69:@2371.4]
  assign _T_4827 = _T_4151 ? 16'h20 : _T_4826; // @[Mux.scala 31:69:@2372.4]
  assign _T_4828 = _T_4148 ? 16'h10 : _T_4827; // @[Mux.scala 31:69:@2373.4]
  assign _T_4829 = _T_4145 ? 16'h8 : _T_4828; // @[Mux.scala 31:69:@2374.4]
  assign _T_4830 = _T_4142 ? 16'h4 : _T_4829; // @[Mux.scala 31:69:@2375.4]
  assign _T_4831 = _T_4139 ? 16'h2 : _T_4830; // @[Mux.scala 31:69:@2376.4]
  assign _T_4832 = _T_4136 ? 16'h1 : _T_4831; // @[Mux.scala 31:69:@2377.4]
  assign _T_4833 = _T_4832[0]; // @[OneHot.scala 66:30:@2378.4]
  assign _T_4834 = _T_4832[1]; // @[OneHot.scala 66:30:@2379.4]
  assign _T_4835 = _T_4832[2]; // @[OneHot.scala 66:30:@2380.4]
  assign _T_4836 = _T_4832[3]; // @[OneHot.scala 66:30:@2381.4]
  assign _T_4837 = _T_4832[4]; // @[OneHot.scala 66:30:@2382.4]
  assign _T_4838 = _T_4832[5]; // @[OneHot.scala 66:30:@2383.4]
  assign _T_4839 = _T_4832[6]; // @[OneHot.scala 66:30:@2384.4]
  assign _T_4840 = _T_4832[7]; // @[OneHot.scala 66:30:@2385.4]
  assign _T_4841 = _T_4832[8]; // @[OneHot.scala 66:30:@2386.4]
  assign _T_4842 = _T_4832[9]; // @[OneHot.scala 66:30:@2387.4]
  assign _T_4843 = _T_4832[10]; // @[OneHot.scala 66:30:@2388.4]
  assign _T_4844 = _T_4832[11]; // @[OneHot.scala 66:30:@2389.4]
  assign _T_4845 = _T_4832[12]; // @[OneHot.scala 66:30:@2390.4]
  assign _T_4846 = _T_4832[13]; // @[OneHot.scala 66:30:@2391.4]
  assign _T_4847 = _T_4832[14]; // @[OneHot.scala 66:30:@2392.4]
  assign _T_4848 = _T_4832[15]; // @[OneHot.scala 66:30:@2393.4]
  assign _T_4889 = _T_4136 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2411.4]
  assign _T_4890 = _T_4133 ? 16'h4000 : _T_4889; // @[Mux.scala 31:69:@2412.4]
  assign _T_4891 = _T_4130 ? 16'h2000 : _T_4890; // @[Mux.scala 31:69:@2413.4]
  assign _T_4892 = _T_4127 ? 16'h1000 : _T_4891; // @[Mux.scala 31:69:@2414.4]
  assign _T_4893 = _T_4124 ? 16'h800 : _T_4892; // @[Mux.scala 31:69:@2415.4]
  assign _T_4894 = _T_4121 ? 16'h400 : _T_4893; // @[Mux.scala 31:69:@2416.4]
  assign _T_4895 = _T_4118 ? 16'h200 : _T_4894; // @[Mux.scala 31:69:@2417.4]
  assign _T_4896 = _T_4115 ? 16'h100 : _T_4895; // @[Mux.scala 31:69:@2418.4]
  assign _T_4897 = _T_4160 ? 16'h80 : _T_4896; // @[Mux.scala 31:69:@2419.4]
  assign _T_4898 = _T_4157 ? 16'h40 : _T_4897; // @[Mux.scala 31:69:@2420.4]
  assign _T_4899 = _T_4154 ? 16'h20 : _T_4898; // @[Mux.scala 31:69:@2421.4]
  assign _T_4900 = _T_4151 ? 16'h10 : _T_4899; // @[Mux.scala 31:69:@2422.4]
  assign _T_4901 = _T_4148 ? 16'h8 : _T_4900; // @[Mux.scala 31:69:@2423.4]
  assign _T_4902 = _T_4145 ? 16'h4 : _T_4901; // @[Mux.scala 31:69:@2424.4]
  assign _T_4903 = _T_4142 ? 16'h2 : _T_4902; // @[Mux.scala 31:69:@2425.4]
  assign _T_4904 = _T_4139 ? 16'h1 : _T_4903; // @[Mux.scala 31:69:@2426.4]
  assign _T_4905 = _T_4904[0]; // @[OneHot.scala 66:30:@2427.4]
  assign _T_4906 = _T_4904[1]; // @[OneHot.scala 66:30:@2428.4]
  assign _T_4907 = _T_4904[2]; // @[OneHot.scala 66:30:@2429.4]
  assign _T_4908 = _T_4904[3]; // @[OneHot.scala 66:30:@2430.4]
  assign _T_4909 = _T_4904[4]; // @[OneHot.scala 66:30:@2431.4]
  assign _T_4910 = _T_4904[5]; // @[OneHot.scala 66:30:@2432.4]
  assign _T_4911 = _T_4904[6]; // @[OneHot.scala 66:30:@2433.4]
  assign _T_4912 = _T_4904[7]; // @[OneHot.scala 66:30:@2434.4]
  assign _T_4913 = _T_4904[8]; // @[OneHot.scala 66:30:@2435.4]
  assign _T_4914 = _T_4904[9]; // @[OneHot.scala 66:30:@2436.4]
  assign _T_4915 = _T_4904[10]; // @[OneHot.scala 66:30:@2437.4]
  assign _T_4916 = _T_4904[11]; // @[OneHot.scala 66:30:@2438.4]
  assign _T_4917 = _T_4904[12]; // @[OneHot.scala 66:30:@2439.4]
  assign _T_4918 = _T_4904[13]; // @[OneHot.scala 66:30:@2440.4]
  assign _T_4919 = _T_4904[14]; // @[OneHot.scala 66:30:@2441.4]
  assign _T_4920 = _T_4904[15]; // @[OneHot.scala 66:30:@2442.4]
  assign _T_4961 = _T_4139 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2460.4]
  assign _T_4962 = _T_4136 ? 16'h4000 : _T_4961; // @[Mux.scala 31:69:@2461.4]
  assign _T_4963 = _T_4133 ? 16'h2000 : _T_4962; // @[Mux.scala 31:69:@2462.4]
  assign _T_4964 = _T_4130 ? 16'h1000 : _T_4963; // @[Mux.scala 31:69:@2463.4]
  assign _T_4965 = _T_4127 ? 16'h800 : _T_4964; // @[Mux.scala 31:69:@2464.4]
  assign _T_4966 = _T_4124 ? 16'h400 : _T_4965; // @[Mux.scala 31:69:@2465.4]
  assign _T_4967 = _T_4121 ? 16'h200 : _T_4966; // @[Mux.scala 31:69:@2466.4]
  assign _T_4968 = _T_4118 ? 16'h100 : _T_4967; // @[Mux.scala 31:69:@2467.4]
  assign _T_4969 = _T_4115 ? 16'h80 : _T_4968; // @[Mux.scala 31:69:@2468.4]
  assign _T_4970 = _T_4160 ? 16'h40 : _T_4969; // @[Mux.scala 31:69:@2469.4]
  assign _T_4971 = _T_4157 ? 16'h20 : _T_4970; // @[Mux.scala 31:69:@2470.4]
  assign _T_4972 = _T_4154 ? 16'h10 : _T_4971; // @[Mux.scala 31:69:@2471.4]
  assign _T_4973 = _T_4151 ? 16'h8 : _T_4972; // @[Mux.scala 31:69:@2472.4]
  assign _T_4974 = _T_4148 ? 16'h4 : _T_4973; // @[Mux.scala 31:69:@2473.4]
  assign _T_4975 = _T_4145 ? 16'h2 : _T_4974; // @[Mux.scala 31:69:@2474.4]
  assign _T_4976 = _T_4142 ? 16'h1 : _T_4975; // @[Mux.scala 31:69:@2475.4]
  assign _T_4977 = _T_4976[0]; // @[OneHot.scala 66:30:@2476.4]
  assign _T_4978 = _T_4976[1]; // @[OneHot.scala 66:30:@2477.4]
  assign _T_4979 = _T_4976[2]; // @[OneHot.scala 66:30:@2478.4]
  assign _T_4980 = _T_4976[3]; // @[OneHot.scala 66:30:@2479.4]
  assign _T_4981 = _T_4976[4]; // @[OneHot.scala 66:30:@2480.4]
  assign _T_4982 = _T_4976[5]; // @[OneHot.scala 66:30:@2481.4]
  assign _T_4983 = _T_4976[6]; // @[OneHot.scala 66:30:@2482.4]
  assign _T_4984 = _T_4976[7]; // @[OneHot.scala 66:30:@2483.4]
  assign _T_4985 = _T_4976[8]; // @[OneHot.scala 66:30:@2484.4]
  assign _T_4986 = _T_4976[9]; // @[OneHot.scala 66:30:@2485.4]
  assign _T_4987 = _T_4976[10]; // @[OneHot.scala 66:30:@2486.4]
  assign _T_4988 = _T_4976[11]; // @[OneHot.scala 66:30:@2487.4]
  assign _T_4989 = _T_4976[12]; // @[OneHot.scala 66:30:@2488.4]
  assign _T_4990 = _T_4976[13]; // @[OneHot.scala 66:30:@2489.4]
  assign _T_4991 = _T_4976[14]; // @[OneHot.scala 66:30:@2490.4]
  assign _T_4992 = _T_4976[15]; // @[OneHot.scala 66:30:@2491.4]
  assign _T_5033 = _T_4142 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2509.4]
  assign _T_5034 = _T_4139 ? 16'h4000 : _T_5033; // @[Mux.scala 31:69:@2510.4]
  assign _T_5035 = _T_4136 ? 16'h2000 : _T_5034; // @[Mux.scala 31:69:@2511.4]
  assign _T_5036 = _T_4133 ? 16'h1000 : _T_5035; // @[Mux.scala 31:69:@2512.4]
  assign _T_5037 = _T_4130 ? 16'h800 : _T_5036; // @[Mux.scala 31:69:@2513.4]
  assign _T_5038 = _T_4127 ? 16'h400 : _T_5037; // @[Mux.scala 31:69:@2514.4]
  assign _T_5039 = _T_4124 ? 16'h200 : _T_5038; // @[Mux.scala 31:69:@2515.4]
  assign _T_5040 = _T_4121 ? 16'h100 : _T_5039; // @[Mux.scala 31:69:@2516.4]
  assign _T_5041 = _T_4118 ? 16'h80 : _T_5040; // @[Mux.scala 31:69:@2517.4]
  assign _T_5042 = _T_4115 ? 16'h40 : _T_5041; // @[Mux.scala 31:69:@2518.4]
  assign _T_5043 = _T_4160 ? 16'h20 : _T_5042; // @[Mux.scala 31:69:@2519.4]
  assign _T_5044 = _T_4157 ? 16'h10 : _T_5043; // @[Mux.scala 31:69:@2520.4]
  assign _T_5045 = _T_4154 ? 16'h8 : _T_5044; // @[Mux.scala 31:69:@2521.4]
  assign _T_5046 = _T_4151 ? 16'h4 : _T_5045; // @[Mux.scala 31:69:@2522.4]
  assign _T_5047 = _T_4148 ? 16'h2 : _T_5046; // @[Mux.scala 31:69:@2523.4]
  assign _T_5048 = _T_4145 ? 16'h1 : _T_5047; // @[Mux.scala 31:69:@2524.4]
  assign _T_5049 = _T_5048[0]; // @[OneHot.scala 66:30:@2525.4]
  assign _T_5050 = _T_5048[1]; // @[OneHot.scala 66:30:@2526.4]
  assign _T_5051 = _T_5048[2]; // @[OneHot.scala 66:30:@2527.4]
  assign _T_5052 = _T_5048[3]; // @[OneHot.scala 66:30:@2528.4]
  assign _T_5053 = _T_5048[4]; // @[OneHot.scala 66:30:@2529.4]
  assign _T_5054 = _T_5048[5]; // @[OneHot.scala 66:30:@2530.4]
  assign _T_5055 = _T_5048[6]; // @[OneHot.scala 66:30:@2531.4]
  assign _T_5056 = _T_5048[7]; // @[OneHot.scala 66:30:@2532.4]
  assign _T_5057 = _T_5048[8]; // @[OneHot.scala 66:30:@2533.4]
  assign _T_5058 = _T_5048[9]; // @[OneHot.scala 66:30:@2534.4]
  assign _T_5059 = _T_5048[10]; // @[OneHot.scala 66:30:@2535.4]
  assign _T_5060 = _T_5048[11]; // @[OneHot.scala 66:30:@2536.4]
  assign _T_5061 = _T_5048[12]; // @[OneHot.scala 66:30:@2537.4]
  assign _T_5062 = _T_5048[13]; // @[OneHot.scala 66:30:@2538.4]
  assign _T_5063 = _T_5048[14]; // @[OneHot.scala 66:30:@2539.4]
  assign _T_5064 = _T_5048[15]; // @[OneHot.scala 66:30:@2540.4]
  assign _T_5105 = _T_4145 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2558.4]
  assign _T_5106 = _T_4142 ? 16'h4000 : _T_5105; // @[Mux.scala 31:69:@2559.4]
  assign _T_5107 = _T_4139 ? 16'h2000 : _T_5106; // @[Mux.scala 31:69:@2560.4]
  assign _T_5108 = _T_4136 ? 16'h1000 : _T_5107; // @[Mux.scala 31:69:@2561.4]
  assign _T_5109 = _T_4133 ? 16'h800 : _T_5108; // @[Mux.scala 31:69:@2562.4]
  assign _T_5110 = _T_4130 ? 16'h400 : _T_5109; // @[Mux.scala 31:69:@2563.4]
  assign _T_5111 = _T_4127 ? 16'h200 : _T_5110; // @[Mux.scala 31:69:@2564.4]
  assign _T_5112 = _T_4124 ? 16'h100 : _T_5111; // @[Mux.scala 31:69:@2565.4]
  assign _T_5113 = _T_4121 ? 16'h80 : _T_5112; // @[Mux.scala 31:69:@2566.4]
  assign _T_5114 = _T_4118 ? 16'h40 : _T_5113; // @[Mux.scala 31:69:@2567.4]
  assign _T_5115 = _T_4115 ? 16'h20 : _T_5114; // @[Mux.scala 31:69:@2568.4]
  assign _T_5116 = _T_4160 ? 16'h10 : _T_5115; // @[Mux.scala 31:69:@2569.4]
  assign _T_5117 = _T_4157 ? 16'h8 : _T_5116; // @[Mux.scala 31:69:@2570.4]
  assign _T_5118 = _T_4154 ? 16'h4 : _T_5117; // @[Mux.scala 31:69:@2571.4]
  assign _T_5119 = _T_4151 ? 16'h2 : _T_5118; // @[Mux.scala 31:69:@2572.4]
  assign _T_5120 = _T_4148 ? 16'h1 : _T_5119; // @[Mux.scala 31:69:@2573.4]
  assign _T_5121 = _T_5120[0]; // @[OneHot.scala 66:30:@2574.4]
  assign _T_5122 = _T_5120[1]; // @[OneHot.scala 66:30:@2575.4]
  assign _T_5123 = _T_5120[2]; // @[OneHot.scala 66:30:@2576.4]
  assign _T_5124 = _T_5120[3]; // @[OneHot.scala 66:30:@2577.4]
  assign _T_5125 = _T_5120[4]; // @[OneHot.scala 66:30:@2578.4]
  assign _T_5126 = _T_5120[5]; // @[OneHot.scala 66:30:@2579.4]
  assign _T_5127 = _T_5120[6]; // @[OneHot.scala 66:30:@2580.4]
  assign _T_5128 = _T_5120[7]; // @[OneHot.scala 66:30:@2581.4]
  assign _T_5129 = _T_5120[8]; // @[OneHot.scala 66:30:@2582.4]
  assign _T_5130 = _T_5120[9]; // @[OneHot.scala 66:30:@2583.4]
  assign _T_5131 = _T_5120[10]; // @[OneHot.scala 66:30:@2584.4]
  assign _T_5132 = _T_5120[11]; // @[OneHot.scala 66:30:@2585.4]
  assign _T_5133 = _T_5120[12]; // @[OneHot.scala 66:30:@2586.4]
  assign _T_5134 = _T_5120[13]; // @[OneHot.scala 66:30:@2587.4]
  assign _T_5135 = _T_5120[14]; // @[OneHot.scala 66:30:@2588.4]
  assign _T_5136 = _T_5120[15]; // @[OneHot.scala 66:30:@2589.4]
  assign _T_5177 = _T_4148 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2607.4]
  assign _T_5178 = _T_4145 ? 16'h4000 : _T_5177; // @[Mux.scala 31:69:@2608.4]
  assign _T_5179 = _T_4142 ? 16'h2000 : _T_5178; // @[Mux.scala 31:69:@2609.4]
  assign _T_5180 = _T_4139 ? 16'h1000 : _T_5179; // @[Mux.scala 31:69:@2610.4]
  assign _T_5181 = _T_4136 ? 16'h800 : _T_5180; // @[Mux.scala 31:69:@2611.4]
  assign _T_5182 = _T_4133 ? 16'h400 : _T_5181; // @[Mux.scala 31:69:@2612.4]
  assign _T_5183 = _T_4130 ? 16'h200 : _T_5182; // @[Mux.scala 31:69:@2613.4]
  assign _T_5184 = _T_4127 ? 16'h100 : _T_5183; // @[Mux.scala 31:69:@2614.4]
  assign _T_5185 = _T_4124 ? 16'h80 : _T_5184; // @[Mux.scala 31:69:@2615.4]
  assign _T_5186 = _T_4121 ? 16'h40 : _T_5185; // @[Mux.scala 31:69:@2616.4]
  assign _T_5187 = _T_4118 ? 16'h20 : _T_5186; // @[Mux.scala 31:69:@2617.4]
  assign _T_5188 = _T_4115 ? 16'h10 : _T_5187; // @[Mux.scala 31:69:@2618.4]
  assign _T_5189 = _T_4160 ? 16'h8 : _T_5188; // @[Mux.scala 31:69:@2619.4]
  assign _T_5190 = _T_4157 ? 16'h4 : _T_5189; // @[Mux.scala 31:69:@2620.4]
  assign _T_5191 = _T_4154 ? 16'h2 : _T_5190; // @[Mux.scala 31:69:@2621.4]
  assign _T_5192 = _T_4151 ? 16'h1 : _T_5191; // @[Mux.scala 31:69:@2622.4]
  assign _T_5193 = _T_5192[0]; // @[OneHot.scala 66:30:@2623.4]
  assign _T_5194 = _T_5192[1]; // @[OneHot.scala 66:30:@2624.4]
  assign _T_5195 = _T_5192[2]; // @[OneHot.scala 66:30:@2625.4]
  assign _T_5196 = _T_5192[3]; // @[OneHot.scala 66:30:@2626.4]
  assign _T_5197 = _T_5192[4]; // @[OneHot.scala 66:30:@2627.4]
  assign _T_5198 = _T_5192[5]; // @[OneHot.scala 66:30:@2628.4]
  assign _T_5199 = _T_5192[6]; // @[OneHot.scala 66:30:@2629.4]
  assign _T_5200 = _T_5192[7]; // @[OneHot.scala 66:30:@2630.4]
  assign _T_5201 = _T_5192[8]; // @[OneHot.scala 66:30:@2631.4]
  assign _T_5202 = _T_5192[9]; // @[OneHot.scala 66:30:@2632.4]
  assign _T_5203 = _T_5192[10]; // @[OneHot.scala 66:30:@2633.4]
  assign _T_5204 = _T_5192[11]; // @[OneHot.scala 66:30:@2634.4]
  assign _T_5205 = _T_5192[12]; // @[OneHot.scala 66:30:@2635.4]
  assign _T_5206 = _T_5192[13]; // @[OneHot.scala 66:30:@2636.4]
  assign _T_5207 = _T_5192[14]; // @[OneHot.scala 66:30:@2637.4]
  assign _T_5208 = _T_5192[15]; // @[OneHot.scala 66:30:@2638.4]
  assign _T_5249 = _T_4151 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2656.4]
  assign _T_5250 = _T_4148 ? 16'h4000 : _T_5249; // @[Mux.scala 31:69:@2657.4]
  assign _T_5251 = _T_4145 ? 16'h2000 : _T_5250; // @[Mux.scala 31:69:@2658.4]
  assign _T_5252 = _T_4142 ? 16'h1000 : _T_5251; // @[Mux.scala 31:69:@2659.4]
  assign _T_5253 = _T_4139 ? 16'h800 : _T_5252; // @[Mux.scala 31:69:@2660.4]
  assign _T_5254 = _T_4136 ? 16'h400 : _T_5253; // @[Mux.scala 31:69:@2661.4]
  assign _T_5255 = _T_4133 ? 16'h200 : _T_5254; // @[Mux.scala 31:69:@2662.4]
  assign _T_5256 = _T_4130 ? 16'h100 : _T_5255; // @[Mux.scala 31:69:@2663.4]
  assign _T_5257 = _T_4127 ? 16'h80 : _T_5256; // @[Mux.scala 31:69:@2664.4]
  assign _T_5258 = _T_4124 ? 16'h40 : _T_5257; // @[Mux.scala 31:69:@2665.4]
  assign _T_5259 = _T_4121 ? 16'h20 : _T_5258; // @[Mux.scala 31:69:@2666.4]
  assign _T_5260 = _T_4118 ? 16'h10 : _T_5259; // @[Mux.scala 31:69:@2667.4]
  assign _T_5261 = _T_4115 ? 16'h8 : _T_5260; // @[Mux.scala 31:69:@2668.4]
  assign _T_5262 = _T_4160 ? 16'h4 : _T_5261; // @[Mux.scala 31:69:@2669.4]
  assign _T_5263 = _T_4157 ? 16'h2 : _T_5262; // @[Mux.scala 31:69:@2670.4]
  assign _T_5264 = _T_4154 ? 16'h1 : _T_5263; // @[Mux.scala 31:69:@2671.4]
  assign _T_5265 = _T_5264[0]; // @[OneHot.scala 66:30:@2672.4]
  assign _T_5266 = _T_5264[1]; // @[OneHot.scala 66:30:@2673.4]
  assign _T_5267 = _T_5264[2]; // @[OneHot.scala 66:30:@2674.4]
  assign _T_5268 = _T_5264[3]; // @[OneHot.scala 66:30:@2675.4]
  assign _T_5269 = _T_5264[4]; // @[OneHot.scala 66:30:@2676.4]
  assign _T_5270 = _T_5264[5]; // @[OneHot.scala 66:30:@2677.4]
  assign _T_5271 = _T_5264[6]; // @[OneHot.scala 66:30:@2678.4]
  assign _T_5272 = _T_5264[7]; // @[OneHot.scala 66:30:@2679.4]
  assign _T_5273 = _T_5264[8]; // @[OneHot.scala 66:30:@2680.4]
  assign _T_5274 = _T_5264[9]; // @[OneHot.scala 66:30:@2681.4]
  assign _T_5275 = _T_5264[10]; // @[OneHot.scala 66:30:@2682.4]
  assign _T_5276 = _T_5264[11]; // @[OneHot.scala 66:30:@2683.4]
  assign _T_5277 = _T_5264[12]; // @[OneHot.scala 66:30:@2684.4]
  assign _T_5278 = _T_5264[13]; // @[OneHot.scala 66:30:@2685.4]
  assign _T_5279 = _T_5264[14]; // @[OneHot.scala 66:30:@2686.4]
  assign _T_5280 = _T_5264[15]; // @[OneHot.scala 66:30:@2687.4]
  assign _T_5321 = _T_4154 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2705.4]
  assign _T_5322 = _T_4151 ? 16'h4000 : _T_5321; // @[Mux.scala 31:69:@2706.4]
  assign _T_5323 = _T_4148 ? 16'h2000 : _T_5322; // @[Mux.scala 31:69:@2707.4]
  assign _T_5324 = _T_4145 ? 16'h1000 : _T_5323; // @[Mux.scala 31:69:@2708.4]
  assign _T_5325 = _T_4142 ? 16'h800 : _T_5324; // @[Mux.scala 31:69:@2709.4]
  assign _T_5326 = _T_4139 ? 16'h400 : _T_5325; // @[Mux.scala 31:69:@2710.4]
  assign _T_5327 = _T_4136 ? 16'h200 : _T_5326; // @[Mux.scala 31:69:@2711.4]
  assign _T_5328 = _T_4133 ? 16'h100 : _T_5327; // @[Mux.scala 31:69:@2712.4]
  assign _T_5329 = _T_4130 ? 16'h80 : _T_5328; // @[Mux.scala 31:69:@2713.4]
  assign _T_5330 = _T_4127 ? 16'h40 : _T_5329; // @[Mux.scala 31:69:@2714.4]
  assign _T_5331 = _T_4124 ? 16'h20 : _T_5330; // @[Mux.scala 31:69:@2715.4]
  assign _T_5332 = _T_4121 ? 16'h10 : _T_5331; // @[Mux.scala 31:69:@2716.4]
  assign _T_5333 = _T_4118 ? 16'h8 : _T_5332; // @[Mux.scala 31:69:@2717.4]
  assign _T_5334 = _T_4115 ? 16'h4 : _T_5333; // @[Mux.scala 31:69:@2718.4]
  assign _T_5335 = _T_4160 ? 16'h2 : _T_5334; // @[Mux.scala 31:69:@2719.4]
  assign _T_5336 = _T_4157 ? 16'h1 : _T_5335; // @[Mux.scala 31:69:@2720.4]
  assign _T_5337 = _T_5336[0]; // @[OneHot.scala 66:30:@2721.4]
  assign _T_5338 = _T_5336[1]; // @[OneHot.scala 66:30:@2722.4]
  assign _T_5339 = _T_5336[2]; // @[OneHot.scala 66:30:@2723.4]
  assign _T_5340 = _T_5336[3]; // @[OneHot.scala 66:30:@2724.4]
  assign _T_5341 = _T_5336[4]; // @[OneHot.scala 66:30:@2725.4]
  assign _T_5342 = _T_5336[5]; // @[OneHot.scala 66:30:@2726.4]
  assign _T_5343 = _T_5336[6]; // @[OneHot.scala 66:30:@2727.4]
  assign _T_5344 = _T_5336[7]; // @[OneHot.scala 66:30:@2728.4]
  assign _T_5345 = _T_5336[8]; // @[OneHot.scala 66:30:@2729.4]
  assign _T_5346 = _T_5336[9]; // @[OneHot.scala 66:30:@2730.4]
  assign _T_5347 = _T_5336[10]; // @[OneHot.scala 66:30:@2731.4]
  assign _T_5348 = _T_5336[11]; // @[OneHot.scala 66:30:@2732.4]
  assign _T_5349 = _T_5336[12]; // @[OneHot.scala 66:30:@2733.4]
  assign _T_5350 = _T_5336[13]; // @[OneHot.scala 66:30:@2734.4]
  assign _T_5351 = _T_5336[14]; // @[OneHot.scala 66:30:@2735.4]
  assign _T_5352 = _T_5336[15]; // @[OneHot.scala 66:30:@2736.4]
  assign _T_5393 = _T_4157 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@2754.4]
  assign _T_5394 = _T_4154 ? 16'h4000 : _T_5393; // @[Mux.scala 31:69:@2755.4]
  assign _T_5395 = _T_4151 ? 16'h2000 : _T_5394; // @[Mux.scala 31:69:@2756.4]
  assign _T_5396 = _T_4148 ? 16'h1000 : _T_5395; // @[Mux.scala 31:69:@2757.4]
  assign _T_5397 = _T_4145 ? 16'h800 : _T_5396; // @[Mux.scala 31:69:@2758.4]
  assign _T_5398 = _T_4142 ? 16'h400 : _T_5397; // @[Mux.scala 31:69:@2759.4]
  assign _T_5399 = _T_4139 ? 16'h200 : _T_5398; // @[Mux.scala 31:69:@2760.4]
  assign _T_5400 = _T_4136 ? 16'h100 : _T_5399; // @[Mux.scala 31:69:@2761.4]
  assign _T_5401 = _T_4133 ? 16'h80 : _T_5400; // @[Mux.scala 31:69:@2762.4]
  assign _T_5402 = _T_4130 ? 16'h40 : _T_5401; // @[Mux.scala 31:69:@2763.4]
  assign _T_5403 = _T_4127 ? 16'h20 : _T_5402; // @[Mux.scala 31:69:@2764.4]
  assign _T_5404 = _T_4124 ? 16'h10 : _T_5403; // @[Mux.scala 31:69:@2765.4]
  assign _T_5405 = _T_4121 ? 16'h8 : _T_5404; // @[Mux.scala 31:69:@2766.4]
  assign _T_5406 = _T_4118 ? 16'h4 : _T_5405; // @[Mux.scala 31:69:@2767.4]
  assign _T_5407 = _T_4115 ? 16'h2 : _T_5406; // @[Mux.scala 31:69:@2768.4]
  assign _T_5408 = _T_4160 ? 16'h1 : _T_5407; // @[Mux.scala 31:69:@2769.4]
  assign _T_5409 = _T_5408[0]; // @[OneHot.scala 66:30:@2770.4]
  assign _T_5410 = _T_5408[1]; // @[OneHot.scala 66:30:@2771.4]
  assign _T_5411 = _T_5408[2]; // @[OneHot.scala 66:30:@2772.4]
  assign _T_5412 = _T_5408[3]; // @[OneHot.scala 66:30:@2773.4]
  assign _T_5413 = _T_5408[4]; // @[OneHot.scala 66:30:@2774.4]
  assign _T_5414 = _T_5408[5]; // @[OneHot.scala 66:30:@2775.4]
  assign _T_5415 = _T_5408[6]; // @[OneHot.scala 66:30:@2776.4]
  assign _T_5416 = _T_5408[7]; // @[OneHot.scala 66:30:@2777.4]
  assign _T_5417 = _T_5408[8]; // @[OneHot.scala 66:30:@2778.4]
  assign _T_5418 = _T_5408[9]; // @[OneHot.scala 66:30:@2779.4]
  assign _T_5419 = _T_5408[10]; // @[OneHot.scala 66:30:@2780.4]
  assign _T_5420 = _T_5408[11]; // @[OneHot.scala 66:30:@2781.4]
  assign _T_5421 = _T_5408[12]; // @[OneHot.scala 66:30:@2782.4]
  assign _T_5422 = _T_5408[13]; // @[OneHot.scala 66:30:@2783.4]
  assign _T_5423 = _T_5408[14]; // @[OneHot.scala 66:30:@2784.4]
  assign _T_5424 = _T_5408[15]; // @[OneHot.scala 66:30:@2785.4]
  assign _T_5489 = {_T_4336,_T_4335,_T_4334,_T_4333,_T_4332,_T_4331,_T_4330,_T_4329}; // @[Mux.scala 19:72:@2809.4]
  assign _T_5497 = {_T_4344,_T_4343,_T_4342,_T_4341,_T_4340,_T_4339,_T_4338,_T_4337,_T_5489}; // @[Mux.scala 19:72:@2817.4]
  assign _T_5499 = _T_4257 ? _T_5497 : 16'h0; // @[Mux.scala 19:72:@2818.4]
  assign _T_5506 = {_T_4407,_T_4406,_T_4405,_T_4404,_T_4403,_T_4402,_T_4401,_T_4416}; // @[Mux.scala 19:72:@2825.4]
  assign _T_5514 = {_T_4415,_T_4414,_T_4413,_T_4412,_T_4411,_T_4410,_T_4409,_T_4408,_T_5506}; // @[Mux.scala 19:72:@2833.4]
  assign _T_5516 = _T_4258 ? _T_5514 : 16'h0; // @[Mux.scala 19:72:@2834.4]
  assign _T_5523 = {_T_4478,_T_4477,_T_4476,_T_4475,_T_4474,_T_4473,_T_4488,_T_4487}; // @[Mux.scala 19:72:@2841.4]
  assign _T_5531 = {_T_4486,_T_4485,_T_4484,_T_4483,_T_4482,_T_4481,_T_4480,_T_4479,_T_5523}; // @[Mux.scala 19:72:@2849.4]
  assign _T_5533 = _T_4259 ? _T_5531 : 16'h0; // @[Mux.scala 19:72:@2850.4]
  assign _T_5540 = {_T_4549,_T_4548,_T_4547,_T_4546,_T_4545,_T_4560,_T_4559,_T_4558}; // @[Mux.scala 19:72:@2857.4]
  assign _T_5548 = {_T_4557,_T_4556,_T_4555,_T_4554,_T_4553,_T_4552,_T_4551,_T_4550,_T_5540}; // @[Mux.scala 19:72:@2865.4]
  assign _T_5550 = _T_4260 ? _T_5548 : 16'h0; // @[Mux.scala 19:72:@2866.4]
  assign _T_5557 = {_T_4620,_T_4619,_T_4618,_T_4617,_T_4632,_T_4631,_T_4630,_T_4629}; // @[Mux.scala 19:72:@2873.4]
  assign _T_5565 = {_T_4628,_T_4627,_T_4626,_T_4625,_T_4624,_T_4623,_T_4622,_T_4621,_T_5557}; // @[Mux.scala 19:72:@2881.4]
  assign _T_5567 = _T_4261 ? _T_5565 : 16'h0; // @[Mux.scala 19:72:@2882.4]
  assign _T_5574 = {_T_4691,_T_4690,_T_4689,_T_4704,_T_4703,_T_4702,_T_4701,_T_4700}; // @[Mux.scala 19:72:@2889.4]
  assign _T_5582 = {_T_4699,_T_4698,_T_4697,_T_4696,_T_4695,_T_4694,_T_4693,_T_4692,_T_5574}; // @[Mux.scala 19:72:@2897.4]
  assign _T_5584 = _T_4262 ? _T_5582 : 16'h0; // @[Mux.scala 19:72:@2898.4]
  assign _T_5591 = {_T_4762,_T_4761,_T_4776,_T_4775,_T_4774,_T_4773,_T_4772,_T_4771}; // @[Mux.scala 19:72:@2905.4]
  assign _T_5599 = {_T_4770,_T_4769,_T_4768,_T_4767,_T_4766,_T_4765,_T_4764,_T_4763,_T_5591}; // @[Mux.scala 19:72:@2913.4]
  assign _T_5601 = _T_4263 ? _T_5599 : 16'h0; // @[Mux.scala 19:72:@2914.4]
  assign _T_5608 = {_T_4833,_T_4848,_T_4847,_T_4846,_T_4845,_T_4844,_T_4843,_T_4842}; // @[Mux.scala 19:72:@2921.4]
  assign _T_5616 = {_T_4841,_T_4840,_T_4839,_T_4838,_T_4837,_T_4836,_T_4835,_T_4834,_T_5608}; // @[Mux.scala 19:72:@2929.4]
  assign _T_5618 = _T_4264 ? _T_5616 : 16'h0; // @[Mux.scala 19:72:@2930.4]
  assign _T_5625 = {_T_4920,_T_4919,_T_4918,_T_4917,_T_4916,_T_4915,_T_4914,_T_4913}; // @[Mux.scala 19:72:@2937.4]
  assign _T_5633 = {_T_4912,_T_4911,_T_4910,_T_4909,_T_4908,_T_4907,_T_4906,_T_4905,_T_5625}; // @[Mux.scala 19:72:@2945.4]
  assign _T_5635 = _T_4265 ? _T_5633 : 16'h0; // @[Mux.scala 19:72:@2946.4]
  assign _T_5642 = {_T_4991,_T_4990,_T_4989,_T_4988,_T_4987,_T_4986,_T_4985,_T_4984}; // @[Mux.scala 19:72:@2953.4]
  assign _T_5650 = {_T_4983,_T_4982,_T_4981,_T_4980,_T_4979,_T_4978,_T_4977,_T_4992,_T_5642}; // @[Mux.scala 19:72:@2961.4]
  assign _T_5652 = _T_4266 ? _T_5650 : 16'h0; // @[Mux.scala 19:72:@2962.4]
  assign _T_5659 = {_T_5062,_T_5061,_T_5060,_T_5059,_T_5058,_T_5057,_T_5056,_T_5055}; // @[Mux.scala 19:72:@2969.4]
  assign _T_5667 = {_T_5054,_T_5053,_T_5052,_T_5051,_T_5050,_T_5049,_T_5064,_T_5063,_T_5659}; // @[Mux.scala 19:72:@2977.4]
  assign _T_5669 = _T_4267 ? _T_5667 : 16'h0; // @[Mux.scala 19:72:@2978.4]
  assign _T_5676 = {_T_5133,_T_5132,_T_5131,_T_5130,_T_5129,_T_5128,_T_5127,_T_5126}; // @[Mux.scala 19:72:@2985.4]
  assign _T_5684 = {_T_5125,_T_5124,_T_5123,_T_5122,_T_5121,_T_5136,_T_5135,_T_5134,_T_5676}; // @[Mux.scala 19:72:@2993.4]
  assign _T_5686 = _T_4268 ? _T_5684 : 16'h0; // @[Mux.scala 19:72:@2994.4]
  assign _T_5693 = {_T_5204,_T_5203,_T_5202,_T_5201,_T_5200,_T_5199,_T_5198,_T_5197}; // @[Mux.scala 19:72:@3001.4]
  assign _T_5701 = {_T_5196,_T_5195,_T_5194,_T_5193,_T_5208,_T_5207,_T_5206,_T_5205,_T_5693}; // @[Mux.scala 19:72:@3009.4]
  assign _T_5703 = _T_4269 ? _T_5701 : 16'h0; // @[Mux.scala 19:72:@3010.4]
  assign _T_5710 = {_T_5275,_T_5274,_T_5273,_T_5272,_T_5271,_T_5270,_T_5269,_T_5268}; // @[Mux.scala 19:72:@3017.4]
  assign _T_5718 = {_T_5267,_T_5266,_T_5265,_T_5280,_T_5279,_T_5278,_T_5277,_T_5276,_T_5710}; // @[Mux.scala 19:72:@3025.4]
  assign _T_5720 = _T_4270 ? _T_5718 : 16'h0; // @[Mux.scala 19:72:@3026.4]
  assign _T_5727 = {_T_5346,_T_5345,_T_5344,_T_5343,_T_5342,_T_5341,_T_5340,_T_5339}; // @[Mux.scala 19:72:@3033.4]
  assign _T_5735 = {_T_5338,_T_5337,_T_5352,_T_5351,_T_5350,_T_5349,_T_5348,_T_5347,_T_5727}; // @[Mux.scala 19:72:@3041.4]
  assign _T_5737 = _T_4271 ? _T_5735 : 16'h0; // @[Mux.scala 19:72:@3042.4]
  assign _T_5744 = {_T_5417,_T_5416,_T_5415,_T_5414,_T_5413,_T_5412,_T_5411,_T_5410}; // @[Mux.scala 19:72:@3049.4]
  assign _T_5752 = {_T_5409,_T_5424,_T_5423,_T_5422,_T_5421,_T_5420,_T_5419,_T_5418,_T_5744}; // @[Mux.scala 19:72:@3057.4]
  assign _T_5754 = _T_4272 ? _T_5752 : 16'h0; // @[Mux.scala 19:72:@3058.4]
  assign _T_5755 = _T_5499 | _T_5516; // @[Mux.scala 19:72:@3059.4]
  assign _T_5756 = _T_5755 | _T_5533; // @[Mux.scala 19:72:@3060.4]
  assign _T_5757 = _T_5756 | _T_5550; // @[Mux.scala 19:72:@3061.4]
  assign _T_5758 = _T_5757 | _T_5567; // @[Mux.scala 19:72:@3062.4]
  assign _T_5759 = _T_5758 | _T_5584; // @[Mux.scala 19:72:@3063.4]
  assign _T_5760 = _T_5759 | _T_5601; // @[Mux.scala 19:72:@3064.4]
  assign _T_5761 = _T_5760 | _T_5618; // @[Mux.scala 19:72:@3065.4]
  assign _T_5762 = _T_5761 | _T_5635; // @[Mux.scala 19:72:@3066.4]
  assign _T_5763 = _T_5762 | _T_5652; // @[Mux.scala 19:72:@3067.4]
  assign _T_5764 = _T_5763 | _T_5669; // @[Mux.scala 19:72:@3068.4]
  assign _T_5765 = _T_5764 | _T_5686; // @[Mux.scala 19:72:@3069.4]
  assign _T_5766 = _T_5765 | _T_5703; // @[Mux.scala 19:72:@3070.4]
  assign _T_5767 = _T_5766 | _T_5720; // @[Mux.scala 19:72:@3071.4]
  assign _T_5768 = _T_5767 | _T_5737; // @[Mux.scala 19:72:@3072.4]
  assign _T_5769 = _T_5768 | _T_5754; // @[Mux.scala 19:72:@3073.4]
  assign inputAddrPriorityPorts_0_0 = _T_5769[0]; // @[Mux.scala 19:72:@3077.4]
  assign inputAddrPriorityPorts_0_1 = _T_5769[1]; // @[Mux.scala 19:72:@3079.4]
  assign inputAddrPriorityPorts_0_2 = _T_5769[2]; // @[Mux.scala 19:72:@3081.4]
  assign inputAddrPriorityPorts_0_3 = _T_5769[3]; // @[Mux.scala 19:72:@3083.4]
  assign inputAddrPriorityPorts_0_4 = _T_5769[4]; // @[Mux.scala 19:72:@3085.4]
  assign inputAddrPriorityPorts_0_5 = _T_5769[5]; // @[Mux.scala 19:72:@3087.4]
  assign inputAddrPriorityPorts_0_6 = _T_5769[6]; // @[Mux.scala 19:72:@3089.4]
  assign inputAddrPriorityPorts_0_7 = _T_5769[7]; // @[Mux.scala 19:72:@3091.4]
  assign inputAddrPriorityPorts_0_8 = _T_5769[8]; // @[Mux.scala 19:72:@3093.4]
  assign inputAddrPriorityPorts_0_9 = _T_5769[9]; // @[Mux.scala 19:72:@3095.4]
  assign inputAddrPriorityPorts_0_10 = _T_5769[10]; // @[Mux.scala 19:72:@3097.4]
  assign inputAddrPriorityPorts_0_11 = _T_5769[11]; // @[Mux.scala 19:72:@3099.4]
  assign inputAddrPriorityPorts_0_12 = _T_5769[12]; // @[Mux.scala 19:72:@3101.4]
  assign inputAddrPriorityPorts_0_13 = _T_5769[13]; // @[Mux.scala 19:72:@3103.4]
  assign inputAddrPriorityPorts_0_14 = _T_5769[14]; // @[Mux.scala 19:72:@3105.4]
  assign inputAddrPriorityPorts_0_15 = _T_5769[15]; // @[Mux.scala 19:72:@3107.4]
  assign _T_5971 = _T_4230 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3161.4]
  assign _T_5972 = _T_4227 ? 16'h4000 : _T_5971; // @[Mux.scala 31:69:@3162.4]
  assign _T_5973 = _T_4224 ? 16'h2000 : _T_5972; // @[Mux.scala 31:69:@3163.4]
  assign _T_5974 = _T_4221 ? 16'h1000 : _T_5973; // @[Mux.scala 31:69:@3164.4]
  assign _T_5975 = _T_4218 ? 16'h800 : _T_5974; // @[Mux.scala 31:69:@3165.4]
  assign _T_5976 = _T_4215 ? 16'h400 : _T_5975; // @[Mux.scala 31:69:@3166.4]
  assign _T_5977 = _T_4212 ? 16'h200 : _T_5976; // @[Mux.scala 31:69:@3167.4]
  assign _T_5978 = _T_4209 ? 16'h100 : _T_5977; // @[Mux.scala 31:69:@3168.4]
  assign _T_5979 = _T_4206 ? 16'h80 : _T_5978; // @[Mux.scala 31:69:@3169.4]
  assign _T_5980 = _T_4203 ? 16'h40 : _T_5979; // @[Mux.scala 31:69:@3170.4]
  assign _T_5981 = _T_4200 ? 16'h20 : _T_5980; // @[Mux.scala 31:69:@3171.4]
  assign _T_5982 = _T_4197 ? 16'h10 : _T_5981; // @[Mux.scala 31:69:@3172.4]
  assign _T_5983 = _T_4194 ? 16'h8 : _T_5982; // @[Mux.scala 31:69:@3173.4]
  assign _T_5984 = _T_4191 ? 16'h4 : _T_5983; // @[Mux.scala 31:69:@3174.4]
  assign _T_5985 = _T_4188 ? 16'h2 : _T_5984; // @[Mux.scala 31:69:@3175.4]
  assign _T_5986 = _T_4185 ? 16'h1 : _T_5985; // @[Mux.scala 31:69:@3176.4]
  assign _T_5987 = _T_5986[0]; // @[OneHot.scala 66:30:@3177.4]
  assign _T_5988 = _T_5986[1]; // @[OneHot.scala 66:30:@3178.4]
  assign _T_5989 = _T_5986[2]; // @[OneHot.scala 66:30:@3179.4]
  assign _T_5990 = _T_5986[3]; // @[OneHot.scala 66:30:@3180.4]
  assign _T_5991 = _T_5986[4]; // @[OneHot.scala 66:30:@3181.4]
  assign _T_5992 = _T_5986[5]; // @[OneHot.scala 66:30:@3182.4]
  assign _T_5993 = _T_5986[6]; // @[OneHot.scala 66:30:@3183.4]
  assign _T_5994 = _T_5986[7]; // @[OneHot.scala 66:30:@3184.4]
  assign _T_5995 = _T_5986[8]; // @[OneHot.scala 66:30:@3185.4]
  assign _T_5996 = _T_5986[9]; // @[OneHot.scala 66:30:@3186.4]
  assign _T_5997 = _T_5986[10]; // @[OneHot.scala 66:30:@3187.4]
  assign _T_5998 = _T_5986[11]; // @[OneHot.scala 66:30:@3188.4]
  assign _T_5999 = _T_5986[12]; // @[OneHot.scala 66:30:@3189.4]
  assign _T_6000 = _T_5986[13]; // @[OneHot.scala 66:30:@3190.4]
  assign _T_6001 = _T_5986[14]; // @[OneHot.scala 66:30:@3191.4]
  assign _T_6002 = _T_5986[15]; // @[OneHot.scala 66:30:@3192.4]
  assign _T_6043 = _T_4185 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3210.4]
  assign _T_6044 = _T_4230 ? 16'h4000 : _T_6043; // @[Mux.scala 31:69:@3211.4]
  assign _T_6045 = _T_4227 ? 16'h2000 : _T_6044; // @[Mux.scala 31:69:@3212.4]
  assign _T_6046 = _T_4224 ? 16'h1000 : _T_6045; // @[Mux.scala 31:69:@3213.4]
  assign _T_6047 = _T_4221 ? 16'h800 : _T_6046; // @[Mux.scala 31:69:@3214.4]
  assign _T_6048 = _T_4218 ? 16'h400 : _T_6047; // @[Mux.scala 31:69:@3215.4]
  assign _T_6049 = _T_4215 ? 16'h200 : _T_6048; // @[Mux.scala 31:69:@3216.4]
  assign _T_6050 = _T_4212 ? 16'h100 : _T_6049; // @[Mux.scala 31:69:@3217.4]
  assign _T_6051 = _T_4209 ? 16'h80 : _T_6050; // @[Mux.scala 31:69:@3218.4]
  assign _T_6052 = _T_4206 ? 16'h40 : _T_6051; // @[Mux.scala 31:69:@3219.4]
  assign _T_6053 = _T_4203 ? 16'h20 : _T_6052; // @[Mux.scala 31:69:@3220.4]
  assign _T_6054 = _T_4200 ? 16'h10 : _T_6053; // @[Mux.scala 31:69:@3221.4]
  assign _T_6055 = _T_4197 ? 16'h8 : _T_6054; // @[Mux.scala 31:69:@3222.4]
  assign _T_6056 = _T_4194 ? 16'h4 : _T_6055; // @[Mux.scala 31:69:@3223.4]
  assign _T_6057 = _T_4191 ? 16'h2 : _T_6056; // @[Mux.scala 31:69:@3224.4]
  assign _T_6058 = _T_4188 ? 16'h1 : _T_6057; // @[Mux.scala 31:69:@3225.4]
  assign _T_6059 = _T_6058[0]; // @[OneHot.scala 66:30:@3226.4]
  assign _T_6060 = _T_6058[1]; // @[OneHot.scala 66:30:@3227.4]
  assign _T_6061 = _T_6058[2]; // @[OneHot.scala 66:30:@3228.4]
  assign _T_6062 = _T_6058[3]; // @[OneHot.scala 66:30:@3229.4]
  assign _T_6063 = _T_6058[4]; // @[OneHot.scala 66:30:@3230.4]
  assign _T_6064 = _T_6058[5]; // @[OneHot.scala 66:30:@3231.4]
  assign _T_6065 = _T_6058[6]; // @[OneHot.scala 66:30:@3232.4]
  assign _T_6066 = _T_6058[7]; // @[OneHot.scala 66:30:@3233.4]
  assign _T_6067 = _T_6058[8]; // @[OneHot.scala 66:30:@3234.4]
  assign _T_6068 = _T_6058[9]; // @[OneHot.scala 66:30:@3235.4]
  assign _T_6069 = _T_6058[10]; // @[OneHot.scala 66:30:@3236.4]
  assign _T_6070 = _T_6058[11]; // @[OneHot.scala 66:30:@3237.4]
  assign _T_6071 = _T_6058[12]; // @[OneHot.scala 66:30:@3238.4]
  assign _T_6072 = _T_6058[13]; // @[OneHot.scala 66:30:@3239.4]
  assign _T_6073 = _T_6058[14]; // @[OneHot.scala 66:30:@3240.4]
  assign _T_6074 = _T_6058[15]; // @[OneHot.scala 66:30:@3241.4]
  assign _T_6115 = _T_4188 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3259.4]
  assign _T_6116 = _T_4185 ? 16'h4000 : _T_6115; // @[Mux.scala 31:69:@3260.4]
  assign _T_6117 = _T_4230 ? 16'h2000 : _T_6116; // @[Mux.scala 31:69:@3261.4]
  assign _T_6118 = _T_4227 ? 16'h1000 : _T_6117; // @[Mux.scala 31:69:@3262.4]
  assign _T_6119 = _T_4224 ? 16'h800 : _T_6118; // @[Mux.scala 31:69:@3263.4]
  assign _T_6120 = _T_4221 ? 16'h400 : _T_6119; // @[Mux.scala 31:69:@3264.4]
  assign _T_6121 = _T_4218 ? 16'h200 : _T_6120; // @[Mux.scala 31:69:@3265.4]
  assign _T_6122 = _T_4215 ? 16'h100 : _T_6121; // @[Mux.scala 31:69:@3266.4]
  assign _T_6123 = _T_4212 ? 16'h80 : _T_6122; // @[Mux.scala 31:69:@3267.4]
  assign _T_6124 = _T_4209 ? 16'h40 : _T_6123; // @[Mux.scala 31:69:@3268.4]
  assign _T_6125 = _T_4206 ? 16'h20 : _T_6124; // @[Mux.scala 31:69:@3269.4]
  assign _T_6126 = _T_4203 ? 16'h10 : _T_6125; // @[Mux.scala 31:69:@3270.4]
  assign _T_6127 = _T_4200 ? 16'h8 : _T_6126; // @[Mux.scala 31:69:@3271.4]
  assign _T_6128 = _T_4197 ? 16'h4 : _T_6127; // @[Mux.scala 31:69:@3272.4]
  assign _T_6129 = _T_4194 ? 16'h2 : _T_6128; // @[Mux.scala 31:69:@3273.4]
  assign _T_6130 = _T_4191 ? 16'h1 : _T_6129; // @[Mux.scala 31:69:@3274.4]
  assign _T_6131 = _T_6130[0]; // @[OneHot.scala 66:30:@3275.4]
  assign _T_6132 = _T_6130[1]; // @[OneHot.scala 66:30:@3276.4]
  assign _T_6133 = _T_6130[2]; // @[OneHot.scala 66:30:@3277.4]
  assign _T_6134 = _T_6130[3]; // @[OneHot.scala 66:30:@3278.4]
  assign _T_6135 = _T_6130[4]; // @[OneHot.scala 66:30:@3279.4]
  assign _T_6136 = _T_6130[5]; // @[OneHot.scala 66:30:@3280.4]
  assign _T_6137 = _T_6130[6]; // @[OneHot.scala 66:30:@3281.4]
  assign _T_6138 = _T_6130[7]; // @[OneHot.scala 66:30:@3282.4]
  assign _T_6139 = _T_6130[8]; // @[OneHot.scala 66:30:@3283.4]
  assign _T_6140 = _T_6130[9]; // @[OneHot.scala 66:30:@3284.4]
  assign _T_6141 = _T_6130[10]; // @[OneHot.scala 66:30:@3285.4]
  assign _T_6142 = _T_6130[11]; // @[OneHot.scala 66:30:@3286.4]
  assign _T_6143 = _T_6130[12]; // @[OneHot.scala 66:30:@3287.4]
  assign _T_6144 = _T_6130[13]; // @[OneHot.scala 66:30:@3288.4]
  assign _T_6145 = _T_6130[14]; // @[OneHot.scala 66:30:@3289.4]
  assign _T_6146 = _T_6130[15]; // @[OneHot.scala 66:30:@3290.4]
  assign _T_6187 = _T_4191 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3308.4]
  assign _T_6188 = _T_4188 ? 16'h4000 : _T_6187; // @[Mux.scala 31:69:@3309.4]
  assign _T_6189 = _T_4185 ? 16'h2000 : _T_6188; // @[Mux.scala 31:69:@3310.4]
  assign _T_6190 = _T_4230 ? 16'h1000 : _T_6189; // @[Mux.scala 31:69:@3311.4]
  assign _T_6191 = _T_4227 ? 16'h800 : _T_6190; // @[Mux.scala 31:69:@3312.4]
  assign _T_6192 = _T_4224 ? 16'h400 : _T_6191; // @[Mux.scala 31:69:@3313.4]
  assign _T_6193 = _T_4221 ? 16'h200 : _T_6192; // @[Mux.scala 31:69:@3314.4]
  assign _T_6194 = _T_4218 ? 16'h100 : _T_6193; // @[Mux.scala 31:69:@3315.4]
  assign _T_6195 = _T_4215 ? 16'h80 : _T_6194; // @[Mux.scala 31:69:@3316.4]
  assign _T_6196 = _T_4212 ? 16'h40 : _T_6195; // @[Mux.scala 31:69:@3317.4]
  assign _T_6197 = _T_4209 ? 16'h20 : _T_6196; // @[Mux.scala 31:69:@3318.4]
  assign _T_6198 = _T_4206 ? 16'h10 : _T_6197; // @[Mux.scala 31:69:@3319.4]
  assign _T_6199 = _T_4203 ? 16'h8 : _T_6198; // @[Mux.scala 31:69:@3320.4]
  assign _T_6200 = _T_4200 ? 16'h4 : _T_6199; // @[Mux.scala 31:69:@3321.4]
  assign _T_6201 = _T_4197 ? 16'h2 : _T_6200; // @[Mux.scala 31:69:@3322.4]
  assign _T_6202 = _T_4194 ? 16'h1 : _T_6201; // @[Mux.scala 31:69:@3323.4]
  assign _T_6203 = _T_6202[0]; // @[OneHot.scala 66:30:@3324.4]
  assign _T_6204 = _T_6202[1]; // @[OneHot.scala 66:30:@3325.4]
  assign _T_6205 = _T_6202[2]; // @[OneHot.scala 66:30:@3326.4]
  assign _T_6206 = _T_6202[3]; // @[OneHot.scala 66:30:@3327.4]
  assign _T_6207 = _T_6202[4]; // @[OneHot.scala 66:30:@3328.4]
  assign _T_6208 = _T_6202[5]; // @[OneHot.scala 66:30:@3329.4]
  assign _T_6209 = _T_6202[6]; // @[OneHot.scala 66:30:@3330.4]
  assign _T_6210 = _T_6202[7]; // @[OneHot.scala 66:30:@3331.4]
  assign _T_6211 = _T_6202[8]; // @[OneHot.scala 66:30:@3332.4]
  assign _T_6212 = _T_6202[9]; // @[OneHot.scala 66:30:@3333.4]
  assign _T_6213 = _T_6202[10]; // @[OneHot.scala 66:30:@3334.4]
  assign _T_6214 = _T_6202[11]; // @[OneHot.scala 66:30:@3335.4]
  assign _T_6215 = _T_6202[12]; // @[OneHot.scala 66:30:@3336.4]
  assign _T_6216 = _T_6202[13]; // @[OneHot.scala 66:30:@3337.4]
  assign _T_6217 = _T_6202[14]; // @[OneHot.scala 66:30:@3338.4]
  assign _T_6218 = _T_6202[15]; // @[OneHot.scala 66:30:@3339.4]
  assign _T_6259 = _T_4194 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3357.4]
  assign _T_6260 = _T_4191 ? 16'h4000 : _T_6259; // @[Mux.scala 31:69:@3358.4]
  assign _T_6261 = _T_4188 ? 16'h2000 : _T_6260; // @[Mux.scala 31:69:@3359.4]
  assign _T_6262 = _T_4185 ? 16'h1000 : _T_6261; // @[Mux.scala 31:69:@3360.4]
  assign _T_6263 = _T_4230 ? 16'h800 : _T_6262; // @[Mux.scala 31:69:@3361.4]
  assign _T_6264 = _T_4227 ? 16'h400 : _T_6263; // @[Mux.scala 31:69:@3362.4]
  assign _T_6265 = _T_4224 ? 16'h200 : _T_6264; // @[Mux.scala 31:69:@3363.4]
  assign _T_6266 = _T_4221 ? 16'h100 : _T_6265; // @[Mux.scala 31:69:@3364.4]
  assign _T_6267 = _T_4218 ? 16'h80 : _T_6266; // @[Mux.scala 31:69:@3365.4]
  assign _T_6268 = _T_4215 ? 16'h40 : _T_6267; // @[Mux.scala 31:69:@3366.4]
  assign _T_6269 = _T_4212 ? 16'h20 : _T_6268; // @[Mux.scala 31:69:@3367.4]
  assign _T_6270 = _T_4209 ? 16'h10 : _T_6269; // @[Mux.scala 31:69:@3368.4]
  assign _T_6271 = _T_4206 ? 16'h8 : _T_6270; // @[Mux.scala 31:69:@3369.4]
  assign _T_6272 = _T_4203 ? 16'h4 : _T_6271; // @[Mux.scala 31:69:@3370.4]
  assign _T_6273 = _T_4200 ? 16'h2 : _T_6272; // @[Mux.scala 31:69:@3371.4]
  assign _T_6274 = _T_4197 ? 16'h1 : _T_6273; // @[Mux.scala 31:69:@3372.4]
  assign _T_6275 = _T_6274[0]; // @[OneHot.scala 66:30:@3373.4]
  assign _T_6276 = _T_6274[1]; // @[OneHot.scala 66:30:@3374.4]
  assign _T_6277 = _T_6274[2]; // @[OneHot.scala 66:30:@3375.4]
  assign _T_6278 = _T_6274[3]; // @[OneHot.scala 66:30:@3376.4]
  assign _T_6279 = _T_6274[4]; // @[OneHot.scala 66:30:@3377.4]
  assign _T_6280 = _T_6274[5]; // @[OneHot.scala 66:30:@3378.4]
  assign _T_6281 = _T_6274[6]; // @[OneHot.scala 66:30:@3379.4]
  assign _T_6282 = _T_6274[7]; // @[OneHot.scala 66:30:@3380.4]
  assign _T_6283 = _T_6274[8]; // @[OneHot.scala 66:30:@3381.4]
  assign _T_6284 = _T_6274[9]; // @[OneHot.scala 66:30:@3382.4]
  assign _T_6285 = _T_6274[10]; // @[OneHot.scala 66:30:@3383.4]
  assign _T_6286 = _T_6274[11]; // @[OneHot.scala 66:30:@3384.4]
  assign _T_6287 = _T_6274[12]; // @[OneHot.scala 66:30:@3385.4]
  assign _T_6288 = _T_6274[13]; // @[OneHot.scala 66:30:@3386.4]
  assign _T_6289 = _T_6274[14]; // @[OneHot.scala 66:30:@3387.4]
  assign _T_6290 = _T_6274[15]; // @[OneHot.scala 66:30:@3388.4]
  assign _T_6331 = _T_4197 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3406.4]
  assign _T_6332 = _T_4194 ? 16'h4000 : _T_6331; // @[Mux.scala 31:69:@3407.4]
  assign _T_6333 = _T_4191 ? 16'h2000 : _T_6332; // @[Mux.scala 31:69:@3408.4]
  assign _T_6334 = _T_4188 ? 16'h1000 : _T_6333; // @[Mux.scala 31:69:@3409.4]
  assign _T_6335 = _T_4185 ? 16'h800 : _T_6334; // @[Mux.scala 31:69:@3410.4]
  assign _T_6336 = _T_4230 ? 16'h400 : _T_6335; // @[Mux.scala 31:69:@3411.4]
  assign _T_6337 = _T_4227 ? 16'h200 : _T_6336; // @[Mux.scala 31:69:@3412.4]
  assign _T_6338 = _T_4224 ? 16'h100 : _T_6337; // @[Mux.scala 31:69:@3413.4]
  assign _T_6339 = _T_4221 ? 16'h80 : _T_6338; // @[Mux.scala 31:69:@3414.4]
  assign _T_6340 = _T_4218 ? 16'h40 : _T_6339; // @[Mux.scala 31:69:@3415.4]
  assign _T_6341 = _T_4215 ? 16'h20 : _T_6340; // @[Mux.scala 31:69:@3416.4]
  assign _T_6342 = _T_4212 ? 16'h10 : _T_6341; // @[Mux.scala 31:69:@3417.4]
  assign _T_6343 = _T_4209 ? 16'h8 : _T_6342; // @[Mux.scala 31:69:@3418.4]
  assign _T_6344 = _T_4206 ? 16'h4 : _T_6343; // @[Mux.scala 31:69:@3419.4]
  assign _T_6345 = _T_4203 ? 16'h2 : _T_6344; // @[Mux.scala 31:69:@3420.4]
  assign _T_6346 = _T_4200 ? 16'h1 : _T_6345; // @[Mux.scala 31:69:@3421.4]
  assign _T_6347 = _T_6346[0]; // @[OneHot.scala 66:30:@3422.4]
  assign _T_6348 = _T_6346[1]; // @[OneHot.scala 66:30:@3423.4]
  assign _T_6349 = _T_6346[2]; // @[OneHot.scala 66:30:@3424.4]
  assign _T_6350 = _T_6346[3]; // @[OneHot.scala 66:30:@3425.4]
  assign _T_6351 = _T_6346[4]; // @[OneHot.scala 66:30:@3426.4]
  assign _T_6352 = _T_6346[5]; // @[OneHot.scala 66:30:@3427.4]
  assign _T_6353 = _T_6346[6]; // @[OneHot.scala 66:30:@3428.4]
  assign _T_6354 = _T_6346[7]; // @[OneHot.scala 66:30:@3429.4]
  assign _T_6355 = _T_6346[8]; // @[OneHot.scala 66:30:@3430.4]
  assign _T_6356 = _T_6346[9]; // @[OneHot.scala 66:30:@3431.4]
  assign _T_6357 = _T_6346[10]; // @[OneHot.scala 66:30:@3432.4]
  assign _T_6358 = _T_6346[11]; // @[OneHot.scala 66:30:@3433.4]
  assign _T_6359 = _T_6346[12]; // @[OneHot.scala 66:30:@3434.4]
  assign _T_6360 = _T_6346[13]; // @[OneHot.scala 66:30:@3435.4]
  assign _T_6361 = _T_6346[14]; // @[OneHot.scala 66:30:@3436.4]
  assign _T_6362 = _T_6346[15]; // @[OneHot.scala 66:30:@3437.4]
  assign _T_6403 = _T_4200 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3455.4]
  assign _T_6404 = _T_4197 ? 16'h4000 : _T_6403; // @[Mux.scala 31:69:@3456.4]
  assign _T_6405 = _T_4194 ? 16'h2000 : _T_6404; // @[Mux.scala 31:69:@3457.4]
  assign _T_6406 = _T_4191 ? 16'h1000 : _T_6405; // @[Mux.scala 31:69:@3458.4]
  assign _T_6407 = _T_4188 ? 16'h800 : _T_6406; // @[Mux.scala 31:69:@3459.4]
  assign _T_6408 = _T_4185 ? 16'h400 : _T_6407; // @[Mux.scala 31:69:@3460.4]
  assign _T_6409 = _T_4230 ? 16'h200 : _T_6408; // @[Mux.scala 31:69:@3461.4]
  assign _T_6410 = _T_4227 ? 16'h100 : _T_6409; // @[Mux.scala 31:69:@3462.4]
  assign _T_6411 = _T_4224 ? 16'h80 : _T_6410; // @[Mux.scala 31:69:@3463.4]
  assign _T_6412 = _T_4221 ? 16'h40 : _T_6411; // @[Mux.scala 31:69:@3464.4]
  assign _T_6413 = _T_4218 ? 16'h20 : _T_6412; // @[Mux.scala 31:69:@3465.4]
  assign _T_6414 = _T_4215 ? 16'h10 : _T_6413; // @[Mux.scala 31:69:@3466.4]
  assign _T_6415 = _T_4212 ? 16'h8 : _T_6414; // @[Mux.scala 31:69:@3467.4]
  assign _T_6416 = _T_4209 ? 16'h4 : _T_6415; // @[Mux.scala 31:69:@3468.4]
  assign _T_6417 = _T_4206 ? 16'h2 : _T_6416; // @[Mux.scala 31:69:@3469.4]
  assign _T_6418 = _T_4203 ? 16'h1 : _T_6417; // @[Mux.scala 31:69:@3470.4]
  assign _T_6419 = _T_6418[0]; // @[OneHot.scala 66:30:@3471.4]
  assign _T_6420 = _T_6418[1]; // @[OneHot.scala 66:30:@3472.4]
  assign _T_6421 = _T_6418[2]; // @[OneHot.scala 66:30:@3473.4]
  assign _T_6422 = _T_6418[3]; // @[OneHot.scala 66:30:@3474.4]
  assign _T_6423 = _T_6418[4]; // @[OneHot.scala 66:30:@3475.4]
  assign _T_6424 = _T_6418[5]; // @[OneHot.scala 66:30:@3476.4]
  assign _T_6425 = _T_6418[6]; // @[OneHot.scala 66:30:@3477.4]
  assign _T_6426 = _T_6418[7]; // @[OneHot.scala 66:30:@3478.4]
  assign _T_6427 = _T_6418[8]; // @[OneHot.scala 66:30:@3479.4]
  assign _T_6428 = _T_6418[9]; // @[OneHot.scala 66:30:@3480.4]
  assign _T_6429 = _T_6418[10]; // @[OneHot.scala 66:30:@3481.4]
  assign _T_6430 = _T_6418[11]; // @[OneHot.scala 66:30:@3482.4]
  assign _T_6431 = _T_6418[12]; // @[OneHot.scala 66:30:@3483.4]
  assign _T_6432 = _T_6418[13]; // @[OneHot.scala 66:30:@3484.4]
  assign _T_6433 = _T_6418[14]; // @[OneHot.scala 66:30:@3485.4]
  assign _T_6434 = _T_6418[15]; // @[OneHot.scala 66:30:@3486.4]
  assign _T_6475 = _T_4203 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3504.4]
  assign _T_6476 = _T_4200 ? 16'h4000 : _T_6475; // @[Mux.scala 31:69:@3505.4]
  assign _T_6477 = _T_4197 ? 16'h2000 : _T_6476; // @[Mux.scala 31:69:@3506.4]
  assign _T_6478 = _T_4194 ? 16'h1000 : _T_6477; // @[Mux.scala 31:69:@3507.4]
  assign _T_6479 = _T_4191 ? 16'h800 : _T_6478; // @[Mux.scala 31:69:@3508.4]
  assign _T_6480 = _T_4188 ? 16'h400 : _T_6479; // @[Mux.scala 31:69:@3509.4]
  assign _T_6481 = _T_4185 ? 16'h200 : _T_6480; // @[Mux.scala 31:69:@3510.4]
  assign _T_6482 = _T_4230 ? 16'h100 : _T_6481; // @[Mux.scala 31:69:@3511.4]
  assign _T_6483 = _T_4227 ? 16'h80 : _T_6482; // @[Mux.scala 31:69:@3512.4]
  assign _T_6484 = _T_4224 ? 16'h40 : _T_6483; // @[Mux.scala 31:69:@3513.4]
  assign _T_6485 = _T_4221 ? 16'h20 : _T_6484; // @[Mux.scala 31:69:@3514.4]
  assign _T_6486 = _T_4218 ? 16'h10 : _T_6485; // @[Mux.scala 31:69:@3515.4]
  assign _T_6487 = _T_4215 ? 16'h8 : _T_6486; // @[Mux.scala 31:69:@3516.4]
  assign _T_6488 = _T_4212 ? 16'h4 : _T_6487; // @[Mux.scala 31:69:@3517.4]
  assign _T_6489 = _T_4209 ? 16'h2 : _T_6488; // @[Mux.scala 31:69:@3518.4]
  assign _T_6490 = _T_4206 ? 16'h1 : _T_6489; // @[Mux.scala 31:69:@3519.4]
  assign _T_6491 = _T_6490[0]; // @[OneHot.scala 66:30:@3520.4]
  assign _T_6492 = _T_6490[1]; // @[OneHot.scala 66:30:@3521.4]
  assign _T_6493 = _T_6490[2]; // @[OneHot.scala 66:30:@3522.4]
  assign _T_6494 = _T_6490[3]; // @[OneHot.scala 66:30:@3523.4]
  assign _T_6495 = _T_6490[4]; // @[OneHot.scala 66:30:@3524.4]
  assign _T_6496 = _T_6490[5]; // @[OneHot.scala 66:30:@3525.4]
  assign _T_6497 = _T_6490[6]; // @[OneHot.scala 66:30:@3526.4]
  assign _T_6498 = _T_6490[7]; // @[OneHot.scala 66:30:@3527.4]
  assign _T_6499 = _T_6490[8]; // @[OneHot.scala 66:30:@3528.4]
  assign _T_6500 = _T_6490[9]; // @[OneHot.scala 66:30:@3529.4]
  assign _T_6501 = _T_6490[10]; // @[OneHot.scala 66:30:@3530.4]
  assign _T_6502 = _T_6490[11]; // @[OneHot.scala 66:30:@3531.4]
  assign _T_6503 = _T_6490[12]; // @[OneHot.scala 66:30:@3532.4]
  assign _T_6504 = _T_6490[13]; // @[OneHot.scala 66:30:@3533.4]
  assign _T_6505 = _T_6490[14]; // @[OneHot.scala 66:30:@3534.4]
  assign _T_6506 = _T_6490[15]; // @[OneHot.scala 66:30:@3535.4]
  assign _T_6547 = _T_4206 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3553.4]
  assign _T_6548 = _T_4203 ? 16'h4000 : _T_6547; // @[Mux.scala 31:69:@3554.4]
  assign _T_6549 = _T_4200 ? 16'h2000 : _T_6548; // @[Mux.scala 31:69:@3555.4]
  assign _T_6550 = _T_4197 ? 16'h1000 : _T_6549; // @[Mux.scala 31:69:@3556.4]
  assign _T_6551 = _T_4194 ? 16'h800 : _T_6550; // @[Mux.scala 31:69:@3557.4]
  assign _T_6552 = _T_4191 ? 16'h400 : _T_6551; // @[Mux.scala 31:69:@3558.4]
  assign _T_6553 = _T_4188 ? 16'h200 : _T_6552; // @[Mux.scala 31:69:@3559.4]
  assign _T_6554 = _T_4185 ? 16'h100 : _T_6553; // @[Mux.scala 31:69:@3560.4]
  assign _T_6555 = _T_4230 ? 16'h80 : _T_6554; // @[Mux.scala 31:69:@3561.4]
  assign _T_6556 = _T_4227 ? 16'h40 : _T_6555; // @[Mux.scala 31:69:@3562.4]
  assign _T_6557 = _T_4224 ? 16'h20 : _T_6556; // @[Mux.scala 31:69:@3563.4]
  assign _T_6558 = _T_4221 ? 16'h10 : _T_6557; // @[Mux.scala 31:69:@3564.4]
  assign _T_6559 = _T_4218 ? 16'h8 : _T_6558; // @[Mux.scala 31:69:@3565.4]
  assign _T_6560 = _T_4215 ? 16'h4 : _T_6559; // @[Mux.scala 31:69:@3566.4]
  assign _T_6561 = _T_4212 ? 16'h2 : _T_6560; // @[Mux.scala 31:69:@3567.4]
  assign _T_6562 = _T_4209 ? 16'h1 : _T_6561; // @[Mux.scala 31:69:@3568.4]
  assign _T_6563 = _T_6562[0]; // @[OneHot.scala 66:30:@3569.4]
  assign _T_6564 = _T_6562[1]; // @[OneHot.scala 66:30:@3570.4]
  assign _T_6565 = _T_6562[2]; // @[OneHot.scala 66:30:@3571.4]
  assign _T_6566 = _T_6562[3]; // @[OneHot.scala 66:30:@3572.4]
  assign _T_6567 = _T_6562[4]; // @[OneHot.scala 66:30:@3573.4]
  assign _T_6568 = _T_6562[5]; // @[OneHot.scala 66:30:@3574.4]
  assign _T_6569 = _T_6562[6]; // @[OneHot.scala 66:30:@3575.4]
  assign _T_6570 = _T_6562[7]; // @[OneHot.scala 66:30:@3576.4]
  assign _T_6571 = _T_6562[8]; // @[OneHot.scala 66:30:@3577.4]
  assign _T_6572 = _T_6562[9]; // @[OneHot.scala 66:30:@3578.4]
  assign _T_6573 = _T_6562[10]; // @[OneHot.scala 66:30:@3579.4]
  assign _T_6574 = _T_6562[11]; // @[OneHot.scala 66:30:@3580.4]
  assign _T_6575 = _T_6562[12]; // @[OneHot.scala 66:30:@3581.4]
  assign _T_6576 = _T_6562[13]; // @[OneHot.scala 66:30:@3582.4]
  assign _T_6577 = _T_6562[14]; // @[OneHot.scala 66:30:@3583.4]
  assign _T_6578 = _T_6562[15]; // @[OneHot.scala 66:30:@3584.4]
  assign _T_6619 = _T_4209 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3602.4]
  assign _T_6620 = _T_4206 ? 16'h4000 : _T_6619; // @[Mux.scala 31:69:@3603.4]
  assign _T_6621 = _T_4203 ? 16'h2000 : _T_6620; // @[Mux.scala 31:69:@3604.4]
  assign _T_6622 = _T_4200 ? 16'h1000 : _T_6621; // @[Mux.scala 31:69:@3605.4]
  assign _T_6623 = _T_4197 ? 16'h800 : _T_6622; // @[Mux.scala 31:69:@3606.4]
  assign _T_6624 = _T_4194 ? 16'h400 : _T_6623; // @[Mux.scala 31:69:@3607.4]
  assign _T_6625 = _T_4191 ? 16'h200 : _T_6624; // @[Mux.scala 31:69:@3608.4]
  assign _T_6626 = _T_4188 ? 16'h100 : _T_6625; // @[Mux.scala 31:69:@3609.4]
  assign _T_6627 = _T_4185 ? 16'h80 : _T_6626; // @[Mux.scala 31:69:@3610.4]
  assign _T_6628 = _T_4230 ? 16'h40 : _T_6627; // @[Mux.scala 31:69:@3611.4]
  assign _T_6629 = _T_4227 ? 16'h20 : _T_6628; // @[Mux.scala 31:69:@3612.4]
  assign _T_6630 = _T_4224 ? 16'h10 : _T_6629; // @[Mux.scala 31:69:@3613.4]
  assign _T_6631 = _T_4221 ? 16'h8 : _T_6630; // @[Mux.scala 31:69:@3614.4]
  assign _T_6632 = _T_4218 ? 16'h4 : _T_6631; // @[Mux.scala 31:69:@3615.4]
  assign _T_6633 = _T_4215 ? 16'h2 : _T_6632; // @[Mux.scala 31:69:@3616.4]
  assign _T_6634 = _T_4212 ? 16'h1 : _T_6633; // @[Mux.scala 31:69:@3617.4]
  assign _T_6635 = _T_6634[0]; // @[OneHot.scala 66:30:@3618.4]
  assign _T_6636 = _T_6634[1]; // @[OneHot.scala 66:30:@3619.4]
  assign _T_6637 = _T_6634[2]; // @[OneHot.scala 66:30:@3620.4]
  assign _T_6638 = _T_6634[3]; // @[OneHot.scala 66:30:@3621.4]
  assign _T_6639 = _T_6634[4]; // @[OneHot.scala 66:30:@3622.4]
  assign _T_6640 = _T_6634[5]; // @[OneHot.scala 66:30:@3623.4]
  assign _T_6641 = _T_6634[6]; // @[OneHot.scala 66:30:@3624.4]
  assign _T_6642 = _T_6634[7]; // @[OneHot.scala 66:30:@3625.4]
  assign _T_6643 = _T_6634[8]; // @[OneHot.scala 66:30:@3626.4]
  assign _T_6644 = _T_6634[9]; // @[OneHot.scala 66:30:@3627.4]
  assign _T_6645 = _T_6634[10]; // @[OneHot.scala 66:30:@3628.4]
  assign _T_6646 = _T_6634[11]; // @[OneHot.scala 66:30:@3629.4]
  assign _T_6647 = _T_6634[12]; // @[OneHot.scala 66:30:@3630.4]
  assign _T_6648 = _T_6634[13]; // @[OneHot.scala 66:30:@3631.4]
  assign _T_6649 = _T_6634[14]; // @[OneHot.scala 66:30:@3632.4]
  assign _T_6650 = _T_6634[15]; // @[OneHot.scala 66:30:@3633.4]
  assign _T_6691 = _T_4212 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3651.4]
  assign _T_6692 = _T_4209 ? 16'h4000 : _T_6691; // @[Mux.scala 31:69:@3652.4]
  assign _T_6693 = _T_4206 ? 16'h2000 : _T_6692; // @[Mux.scala 31:69:@3653.4]
  assign _T_6694 = _T_4203 ? 16'h1000 : _T_6693; // @[Mux.scala 31:69:@3654.4]
  assign _T_6695 = _T_4200 ? 16'h800 : _T_6694; // @[Mux.scala 31:69:@3655.4]
  assign _T_6696 = _T_4197 ? 16'h400 : _T_6695; // @[Mux.scala 31:69:@3656.4]
  assign _T_6697 = _T_4194 ? 16'h200 : _T_6696; // @[Mux.scala 31:69:@3657.4]
  assign _T_6698 = _T_4191 ? 16'h100 : _T_6697; // @[Mux.scala 31:69:@3658.4]
  assign _T_6699 = _T_4188 ? 16'h80 : _T_6698; // @[Mux.scala 31:69:@3659.4]
  assign _T_6700 = _T_4185 ? 16'h40 : _T_6699; // @[Mux.scala 31:69:@3660.4]
  assign _T_6701 = _T_4230 ? 16'h20 : _T_6700; // @[Mux.scala 31:69:@3661.4]
  assign _T_6702 = _T_4227 ? 16'h10 : _T_6701; // @[Mux.scala 31:69:@3662.4]
  assign _T_6703 = _T_4224 ? 16'h8 : _T_6702; // @[Mux.scala 31:69:@3663.4]
  assign _T_6704 = _T_4221 ? 16'h4 : _T_6703; // @[Mux.scala 31:69:@3664.4]
  assign _T_6705 = _T_4218 ? 16'h2 : _T_6704; // @[Mux.scala 31:69:@3665.4]
  assign _T_6706 = _T_4215 ? 16'h1 : _T_6705; // @[Mux.scala 31:69:@3666.4]
  assign _T_6707 = _T_6706[0]; // @[OneHot.scala 66:30:@3667.4]
  assign _T_6708 = _T_6706[1]; // @[OneHot.scala 66:30:@3668.4]
  assign _T_6709 = _T_6706[2]; // @[OneHot.scala 66:30:@3669.4]
  assign _T_6710 = _T_6706[3]; // @[OneHot.scala 66:30:@3670.4]
  assign _T_6711 = _T_6706[4]; // @[OneHot.scala 66:30:@3671.4]
  assign _T_6712 = _T_6706[5]; // @[OneHot.scala 66:30:@3672.4]
  assign _T_6713 = _T_6706[6]; // @[OneHot.scala 66:30:@3673.4]
  assign _T_6714 = _T_6706[7]; // @[OneHot.scala 66:30:@3674.4]
  assign _T_6715 = _T_6706[8]; // @[OneHot.scala 66:30:@3675.4]
  assign _T_6716 = _T_6706[9]; // @[OneHot.scala 66:30:@3676.4]
  assign _T_6717 = _T_6706[10]; // @[OneHot.scala 66:30:@3677.4]
  assign _T_6718 = _T_6706[11]; // @[OneHot.scala 66:30:@3678.4]
  assign _T_6719 = _T_6706[12]; // @[OneHot.scala 66:30:@3679.4]
  assign _T_6720 = _T_6706[13]; // @[OneHot.scala 66:30:@3680.4]
  assign _T_6721 = _T_6706[14]; // @[OneHot.scala 66:30:@3681.4]
  assign _T_6722 = _T_6706[15]; // @[OneHot.scala 66:30:@3682.4]
  assign _T_6763 = _T_4215 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3700.4]
  assign _T_6764 = _T_4212 ? 16'h4000 : _T_6763; // @[Mux.scala 31:69:@3701.4]
  assign _T_6765 = _T_4209 ? 16'h2000 : _T_6764; // @[Mux.scala 31:69:@3702.4]
  assign _T_6766 = _T_4206 ? 16'h1000 : _T_6765; // @[Mux.scala 31:69:@3703.4]
  assign _T_6767 = _T_4203 ? 16'h800 : _T_6766; // @[Mux.scala 31:69:@3704.4]
  assign _T_6768 = _T_4200 ? 16'h400 : _T_6767; // @[Mux.scala 31:69:@3705.4]
  assign _T_6769 = _T_4197 ? 16'h200 : _T_6768; // @[Mux.scala 31:69:@3706.4]
  assign _T_6770 = _T_4194 ? 16'h100 : _T_6769; // @[Mux.scala 31:69:@3707.4]
  assign _T_6771 = _T_4191 ? 16'h80 : _T_6770; // @[Mux.scala 31:69:@3708.4]
  assign _T_6772 = _T_4188 ? 16'h40 : _T_6771; // @[Mux.scala 31:69:@3709.4]
  assign _T_6773 = _T_4185 ? 16'h20 : _T_6772; // @[Mux.scala 31:69:@3710.4]
  assign _T_6774 = _T_4230 ? 16'h10 : _T_6773; // @[Mux.scala 31:69:@3711.4]
  assign _T_6775 = _T_4227 ? 16'h8 : _T_6774; // @[Mux.scala 31:69:@3712.4]
  assign _T_6776 = _T_4224 ? 16'h4 : _T_6775; // @[Mux.scala 31:69:@3713.4]
  assign _T_6777 = _T_4221 ? 16'h2 : _T_6776; // @[Mux.scala 31:69:@3714.4]
  assign _T_6778 = _T_4218 ? 16'h1 : _T_6777; // @[Mux.scala 31:69:@3715.4]
  assign _T_6779 = _T_6778[0]; // @[OneHot.scala 66:30:@3716.4]
  assign _T_6780 = _T_6778[1]; // @[OneHot.scala 66:30:@3717.4]
  assign _T_6781 = _T_6778[2]; // @[OneHot.scala 66:30:@3718.4]
  assign _T_6782 = _T_6778[3]; // @[OneHot.scala 66:30:@3719.4]
  assign _T_6783 = _T_6778[4]; // @[OneHot.scala 66:30:@3720.4]
  assign _T_6784 = _T_6778[5]; // @[OneHot.scala 66:30:@3721.4]
  assign _T_6785 = _T_6778[6]; // @[OneHot.scala 66:30:@3722.4]
  assign _T_6786 = _T_6778[7]; // @[OneHot.scala 66:30:@3723.4]
  assign _T_6787 = _T_6778[8]; // @[OneHot.scala 66:30:@3724.4]
  assign _T_6788 = _T_6778[9]; // @[OneHot.scala 66:30:@3725.4]
  assign _T_6789 = _T_6778[10]; // @[OneHot.scala 66:30:@3726.4]
  assign _T_6790 = _T_6778[11]; // @[OneHot.scala 66:30:@3727.4]
  assign _T_6791 = _T_6778[12]; // @[OneHot.scala 66:30:@3728.4]
  assign _T_6792 = _T_6778[13]; // @[OneHot.scala 66:30:@3729.4]
  assign _T_6793 = _T_6778[14]; // @[OneHot.scala 66:30:@3730.4]
  assign _T_6794 = _T_6778[15]; // @[OneHot.scala 66:30:@3731.4]
  assign _T_6835 = _T_4218 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3749.4]
  assign _T_6836 = _T_4215 ? 16'h4000 : _T_6835; // @[Mux.scala 31:69:@3750.4]
  assign _T_6837 = _T_4212 ? 16'h2000 : _T_6836; // @[Mux.scala 31:69:@3751.4]
  assign _T_6838 = _T_4209 ? 16'h1000 : _T_6837; // @[Mux.scala 31:69:@3752.4]
  assign _T_6839 = _T_4206 ? 16'h800 : _T_6838; // @[Mux.scala 31:69:@3753.4]
  assign _T_6840 = _T_4203 ? 16'h400 : _T_6839; // @[Mux.scala 31:69:@3754.4]
  assign _T_6841 = _T_4200 ? 16'h200 : _T_6840; // @[Mux.scala 31:69:@3755.4]
  assign _T_6842 = _T_4197 ? 16'h100 : _T_6841; // @[Mux.scala 31:69:@3756.4]
  assign _T_6843 = _T_4194 ? 16'h80 : _T_6842; // @[Mux.scala 31:69:@3757.4]
  assign _T_6844 = _T_4191 ? 16'h40 : _T_6843; // @[Mux.scala 31:69:@3758.4]
  assign _T_6845 = _T_4188 ? 16'h20 : _T_6844; // @[Mux.scala 31:69:@3759.4]
  assign _T_6846 = _T_4185 ? 16'h10 : _T_6845; // @[Mux.scala 31:69:@3760.4]
  assign _T_6847 = _T_4230 ? 16'h8 : _T_6846; // @[Mux.scala 31:69:@3761.4]
  assign _T_6848 = _T_4227 ? 16'h4 : _T_6847; // @[Mux.scala 31:69:@3762.4]
  assign _T_6849 = _T_4224 ? 16'h2 : _T_6848; // @[Mux.scala 31:69:@3763.4]
  assign _T_6850 = _T_4221 ? 16'h1 : _T_6849; // @[Mux.scala 31:69:@3764.4]
  assign _T_6851 = _T_6850[0]; // @[OneHot.scala 66:30:@3765.4]
  assign _T_6852 = _T_6850[1]; // @[OneHot.scala 66:30:@3766.4]
  assign _T_6853 = _T_6850[2]; // @[OneHot.scala 66:30:@3767.4]
  assign _T_6854 = _T_6850[3]; // @[OneHot.scala 66:30:@3768.4]
  assign _T_6855 = _T_6850[4]; // @[OneHot.scala 66:30:@3769.4]
  assign _T_6856 = _T_6850[5]; // @[OneHot.scala 66:30:@3770.4]
  assign _T_6857 = _T_6850[6]; // @[OneHot.scala 66:30:@3771.4]
  assign _T_6858 = _T_6850[7]; // @[OneHot.scala 66:30:@3772.4]
  assign _T_6859 = _T_6850[8]; // @[OneHot.scala 66:30:@3773.4]
  assign _T_6860 = _T_6850[9]; // @[OneHot.scala 66:30:@3774.4]
  assign _T_6861 = _T_6850[10]; // @[OneHot.scala 66:30:@3775.4]
  assign _T_6862 = _T_6850[11]; // @[OneHot.scala 66:30:@3776.4]
  assign _T_6863 = _T_6850[12]; // @[OneHot.scala 66:30:@3777.4]
  assign _T_6864 = _T_6850[13]; // @[OneHot.scala 66:30:@3778.4]
  assign _T_6865 = _T_6850[14]; // @[OneHot.scala 66:30:@3779.4]
  assign _T_6866 = _T_6850[15]; // @[OneHot.scala 66:30:@3780.4]
  assign _T_6907 = _T_4221 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3798.4]
  assign _T_6908 = _T_4218 ? 16'h4000 : _T_6907; // @[Mux.scala 31:69:@3799.4]
  assign _T_6909 = _T_4215 ? 16'h2000 : _T_6908; // @[Mux.scala 31:69:@3800.4]
  assign _T_6910 = _T_4212 ? 16'h1000 : _T_6909; // @[Mux.scala 31:69:@3801.4]
  assign _T_6911 = _T_4209 ? 16'h800 : _T_6910; // @[Mux.scala 31:69:@3802.4]
  assign _T_6912 = _T_4206 ? 16'h400 : _T_6911; // @[Mux.scala 31:69:@3803.4]
  assign _T_6913 = _T_4203 ? 16'h200 : _T_6912; // @[Mux.scala 31:69:@3804.4]
  assign _T_6914 = _T_4200 ? 16'h100 : _T_6913; // @[Mux.scala 31:69:@3805.4]
  assign _T_6915 = _T_4197 ? 16'h80 : _T_6914; // @[Mux.scala 31:69:@3806.4]
  assign _T_6916 = _T_4194 ? 16'h40 : _T_6915; // @[Mux.scala 31:69:@3807.4]
  assign _T_6917 = _T_4191 ? 16'h20 : _T_6916; // @[Mux.scala 31:69:@3808.4]
  assign _T_6918 = _T_4188 ? 16'h10 : _T_6917; // @[Mux.scala 31:69:@3809.4]
  assign _T_6919 = _T_4185 ? 16'h8 : _T_6918; // @[Mux.scala 31:69:@3810.4]
  assign _T_6920 = _T_4230 ? 16'h4 : _T_6919; // @[Mux.scala 31:69:@3811.4]
  assign _T_6921 = _T_4227 ? 16'h2 : _T_6920; // @[Mux.scala 31:69:@3812.4]
  assign _T_6922 = _T_4224 ? 16'h1 : _T_6921; // @[Mux.scala 31:69:@3813.4]
  assign _T_6923 = _T_6922[0]; // @[OneHot.scala 66:30:@3814.4]
  assign _T_6924 = _T_6922[1]; // @[OneHot.scala 66:30:@3815.4]
  assign _T_6925 = _T_6922[2]; // @[OneHot.scala 66:30:@3816.4]
  assign _T_6926 = _T_6922[3]; // @[OneHot.scala 66:30:@3817.4]
  assign _T_6927 = _T_6922[4]; // @[OneHot.scala 66:30:@3818.4]
  assign _T_6928 = _T_6922[5]; // @[OneHot.scala 66:30:@3819.4]
  assign _T_6929 = _T_6922[6]; // @[OneHot.scala 66:30:@3820.4]
  assign _T_6930 = _T_6922[7]; // @[OneHot.scala 66:30:@3821.4]
  assign _T_6931 = _T_6922[8]; // @[OneHot.scala 66:30:@3822.4]
  assign _T_6932 = _T_6922[9]; // @[OneHot.scala 66:30:@3823.4]
  assign _T_6933 = _T_6922[10]; // @[OneHot.scala 66:30:@3824.4]
  assign _T_6934 = _T_6922[11]; // @[OneHot.scala 66:30:@3825.4]
  assign _T_6935 = _T_6922[12]; // @[OneHot.scala 66:30:@3826.4]
  assign _T_6936 = _T_6922[13]; // @[OneHot.scala 66:30:@3827.4]
  assign _T_6937 = _T_6922[14]; // @[OneHot.scala 66:30:@3828.4]
  assign _T_6938 = _T_6922[15]; // @[OneHot.scala 66:30:@3829.4]
  assign _T_6979 = _T_4224 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3847.4]
  assign _T_6980 = _T_4221 ? 16'h4000 : _T_6979; // @[Mux.scala 31:69:@3848.4]
  assign _T_6981 = _T_4218 ? 16'h2000 : _T_6980; // @[Mux.scala 31:69:@3849.4]
  assign _T_6982 = _T_4215 ? 16'h1000 : _T_6981; // @[Mux.scala 31:69:@3850.4]
  assign _T_6983 = _T_4212 ? 16'h800 : _T_6982; // @[Mux.scala 31:69:@3851.4]
  assign _T_6984 = _T_4209 ? 16'h400 : _T_6983; // @[Mux.scala 31:69:@3852.4]
  assign _T_6985 = _T_4206 ? 16'h200 : _T_6984; // @[Mux.scala 31:69:@3853.4]
  assign _T_6986 = _T_4203 ? 16'h100 : _T_6985; // @[Mux.scala 31:69:@3854.4]
  assign _T_6987 = _T_4200 ? 16'h80 : _T_6986; // @[Mux.scala 31:69:@3855.4]
  assign _T_6988 = _T_4197 ? 16'h40 : _T_6987; // @[Mux.scala 31:69:@3856.4]
  assign _T_6989 = _T_4194 ? 16'h20 : _T_6988; // @[Mux.scala 31:69:@3857.4]
  assign _T_6990 = _T_4191 ? 16'h10 : _T_6989; // @[Mux.scala 31:69:@3858.4]
  assign _T_6991 = _T_4188 ? 16'h8 : _T_6990; // @[Mux.scala 31:69:@3859.4]
  assign _T_6992 = _T_4185 ? 16'h4 : _T_6991; // @[Mux.scala 31:69:@3860.4]
  assign _T_6993 = _T_4230 ? 16'h2 : _T_6992; // @[Mux.scala 31:69:@3861.4]
  assign _T_6994 = _T_4227 ? 16'h1 : _T_6993; // @[Mux.scala 31:69:@3862.4]
  assign _T_6995 = _T_6994[0]; // @[OneHot.scala 66:30:@3863.4]
  assign _T_6996 = _T_6994[1]; // @[OneHot.scala 66:30:@3864.4]
  assign _T_6997 = _T_6994[2]; // @[OneHot.scala 66:30:@3865.4]
  assign _T_6998 = _T_6994[3]; // @[OneHot.scala 66:30:@3866.4]
  assign _T_6999 = _T_6994[4]; // @[OneHot.scala 66:30:@3867.4]
  assign _T_7000 = _T_6994[5]; // @[OneHot.scala 66:30:@3868.4]
  assign _T_7001 = _T_6994[6]; // @[OneHot.scala 66:30:@3869.4]
  assign _T_7002 = _T_6994[7]; // @[OneHot.scala 66:30:@3870.4]
  assign _T_7003 = _T_6994[8]; // @[OneHot.scala 66:30:@3871.4]
  assign _T_7004 = _T_6994[9]; // @[OneHot.scala 66:30:@3872.4]
  assign _T_7005 = _T_6994[10]; // @[OneHot.scala 66:30:@3873.4]
  assign _T_7006 = _T_6994[11]; // @[OneHot.scala 66:30:@3874.4]
  assign _T_7007 = _T_6994[12]; // @[OneHot.scala 66:30:@3875.4]
  assign _T_7008 = _T_6994[13]; // @[OneHot.scala 66:30:@3876.4]
  assign _T_7009 = _T_6994[14]; // @[OneHot.scala 66:30:@3877.4]
  assign _T_7010 = _T_6994[15]; // @[OneHot.scala 66:30:@3878.4]
  assign _T_7051 = _T_4227 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@3896.4]
  assign _T_7052 = _T_4224 ? 16'h4000 : _T_7051; // @[Mux.scala 31:69:@3897.4]
  assign _T_7053 = _T_4221 ? 16'h2000 : _T_7052; // @[Mux.scala 31:69:@3898.4]
  assign _T_7054 = _T_4218 ? 16'h1000 : _T_7053; // @[Mux.scala 31:69:@3899.4]
  assign _T_7055 = _T_4215 ? 16'h800 : _T_7054; // @[Mux.scala 31:69:@3900.4]
  assign _T_7056 = _T_4212 ? 16'h400 : _T_7055; // @[Mux.scala 31:69:@3901.4]
  assign _T_7057 = _T_4209 ? 16'h200 : _T_7056; // @[Mux.scala 31:69:@3902.4]
  assign _T_7058 = _T_4206 ? 16'h100 : _T_7057; // @[Mux.scala 31:69:@3903.4]
  assign _T_7059 = _T_4203 ? 16'h80 : _T_7058; // @[Mux.scala 31:69:@3904.4]
  assign _T_7060 = _T_4200 ? 16'h40 : _T_7059; // @[Mux.scala 31:69:@3905.4]
  assign _T_7061 = _T_4197 ? 16'h20 : _T_7060; // @[Mux.scala 31:69:@3906.4]
  assign _T_7062 = _T_4194 ? 16'h10 : _T_7061; // @[Mux.scala 31:69:@3907.4]
  assign _T_7063 = _T_4191 ? 16'h8 : _T_7062; // @[Mux.scala 31:69:@3908.4]
  assign _T_7064 = _T_4188 ? 16'h4 : _T_7063; // @[Mux.scala 31:69:@3909.4]
  assign _T_7065 = _T_4185 ? 16'h2 : _T_7064; // @[Mux.scala 31:69:@3910.4]
  assign _T_7066 = _T_4230 ? 16'h1 : _T_7065; // @[Mux.scala 31:69:@3911.4]
  assign _T_7067 = _T_7066[0]; // @[OneHot.scala 66:30:@3912.4]
  assign _T_7068 = _T_7066[1]; // @[OneHot.scala 66:30:@3913.4]
  assign _T_7069 = _T_7066[2]; // @[OneHot.scala 66:30:@3914.4]
  assign _T_7070 = _T_7066[3]; // @[OneHot.scala 66:30:@3915.4]
  assign _T_7071 = _T_7066[4]; // @[OneHot.scala 66:30:@3916.4]
  assign _T_7072 = _T_7066[5]; // @[OneHot.scala 66:30:@3917.4]
  assign _T_7073 = _T_7066[6]; // @[OneHot.scala 66:30:@3918.4]
  assign _T_7074 = _T_7066[7]; // @[OneHot.scala 66:30:@3919.4]
  assign _T_7075 = _T_7066[8]; // @[OneHot.scala 66:30:@3920.4]
  assign _T_7076 = _T_7066[9]; // @[OneHot.scala 66:30:@3921.4]
  assign _T_7077 = _T_7066[10]; // @[OneHot.scala 66:30:@3922.4]
  assign _T_7078 = _T_7066[11]; // @[OneHot.scala 66:30:@3923.4]
  assign _T_7079 = _T_7066[12]; // @[OneHot.scala 66:30:@3924.4]
  assign _T_7080 = _T_7066[13]; // @[OneHot.scala 66:30:@3925.4]
  assign _T_7081 = _T_7066[14]; // @[OneHot.scala 66:30:@3926.4]
  assign _T_7082 = _T_7066[15]; // @[OneHot.scala 66:30:@3927.4]
  assign _T_7147 = {_T_5994,_T_5993,_T_5992,_T_5991,_T_5990,_T_5989,_T_5988,_T_5987}; // @[Mux.scala 19:72:@3951.4]
  assign _T_7155 = {_T_6002,_T_6001,_T_6000,_T_5999,_T_5998,_T_5997,_T_5996,_T_5995,_T_7147}; // @[Mux.scala 19:72:@3959.4]
  assign _T_7157 = _T_4257 ? _T_7155 : 16'h0; // @[Mux.scala 19:72:@3960.4]
  assign _T_7164 = {_T_6065,_T_6064,_T_6063,_T_6062,_T_6061,_T_6060,_T_6059,_T_6074}; // @[Mux.scala 19:72:@3967.4]
  assign _T_7172 = {_T_6073,_T_6072,_T_6071,_T_6070,_T_6069,_T_6068,_T_6067,_T_6066,_T_7164}; // @[Mux.scala 19:72:@3975.4]
  assign _T_7174 = _T_4258 ? _T_7172 : 16'h0; // @[Mux.scala 19:72:@3976.4]
  assign _T_7181 = {_T_6136,_T_6135,_T_6134,_T_6133,_T_6132,_T_6131,_T_6146,_T_6145}; // @[Mux.scala 19:72:@3983.4]
  assign _T_7189 = {_T_6144,_T_6143,_T_6142,_T_6141,_T_6140,_T_6139,_T_6138,_T_6137,_T_7181}; // @[Mux.scala 19:72:@3991.4]
  assign _T_7191 = _T_4259 ? _T_7189 : 16'h0; // @[Mux.scala 19:72:@3992.4]
  assign _T_7198 = {_T_6207,_T_6206,_T_6205,_T_6204,_T_6203,_T_6218,_T_6217,_T_6216}; // @[Mux.scala 19:72:@3999.4]
  assign _T_7206 = {_T_6215,_T_6214,_T_6213,_T_6212,_T_6211,_T_6210,_T_6209,_T_6208,_T_7198}; // @[Mux.scala 19:72:@4007.4]
  assign _T_7208 = _T_4260 ? _T_7206 : 16'h0; // @[Mux.scala 19:72:@4008.4]
  assign _T_7215 = {_T_6278,_T_6277,_T_6276,_T_6275,_T_6290,_T_6289,_T_6288,_T_6287}; // @[Mux.scala 19:72:@4015.4]
  assign _T_7223 = {_T_6286,_T_6285,_T_6284,_T_6283,_T_6282,_T_6281,_T_6280,_T_6279,_T_7215}; // @[Mux.scala 19:72:@4023.4]
  assign _T_7225 = _T_4261 ? _T_7223 : 16'h0; // @[Mux.scala 19:72:@4024.4]
  assign _T_7232 = {_T_6349,_T_6348,_T_6347,_T_6362,_T_6361,_T_6360,_T_6359,_T_6358}; // @[Mux.scala 19:72:@4031.4]
  assign _T_7240 = {_T_6357,_T_6356,_T_6355,_T_6354,_T_6353,_T_6352,_T_6351,_T_6350,_T_7232}; // @[Mux.scala 19:72:@4039.4]
  assign _T_7242 = _T_4262 ? _T_7240 : 16'h0; // @[Mux.scala 19:72:@4040.4]
  assign _T_7249 = {_T_6420,_T_6419,_T_6434,_T_6433,_T_6432,_T_6431,_T_6430,_T_6429}; // @[Mux.scala 19:72:@4047.4]
  assign _T_7257 = {_T_6428,_T_6427,_T_6426,_T_6425,_T_6424,_T_6423,_T_6422,_T_6421,_T_7249}; // @[Mux.scala 19:72:@4055.4]
  assign _T_7259 = _T_4263 ? _T_7257 : 16'h0; // @[Mux.scala 19:72:@4056.4]
  assign _T_7266 = {_T_6491,_T_6506,_T_6505,_T_6504,_T_6503,_T_6502,_T_6501,_T_6500}; // @[Mux.scala 19:72:@4063.4]
  assign _T_7274 = {_T_6499,_T_6498,_T_6497,_T_6496,_T_6495,_T_6494,_T_6493,_T_6492,_T_7266}; // @[Mux.scala 19:72:@4071.4]
  assign _T_7276 = _T_4264 ? _T_7274 : 16'h0; // @[Mux.scala 19:72:@4072.4]
  assign _T_7283 = {_T_6578,_T_6577,_T_6576,_T_6575,_T_6574,_T_6573,_T_6572,_T_6571}; // @[Mux.scala 19:72:@4079.4]
  assign _T_7291 = {_T_6570,_T_6569,_T_6568,_T_6567,_T_6566,_T_6565,_T_6564,_T_6563,_T_7283}; // @[Mux.scala 19:72:@4087.4]
  assign _T_7293 = _T_4265 ? _T_7291 : 16'h0; // @[Mux.scala 19:72:@4088.4]
  assign _T_7300 = {_T_6649,_T_6648,_T_6647,_T_6646,_T_6645,_T_6644,_T_6643,_T_6642}; // @[Mux.scala 19:72:@4095.4]
  assign _T_7308 = {_T_6641,_T_6640,_T_6639,_T_6638,_T_6637,_T_6636,_T_6635,_T_6650,_T_7300}; // @[Mux.scala 19:72:@4103.4]
  assign _T_7310 = _T_4266 ? _T_7308 : 16'h0; // @[Mux.scala 19:72:@4104.4]
  assign _T_7317 = {_T_6720,_T_6719,_T_6718,_T_6717,_T_6716,_T_6715,_T_6714,_T_6713}; // @[Mux.scala 19:72:@4111.4]
  assign _T_7325 = {_T_6712,_T_6711,_T_6710,_T_6709,_T_6708,_T_6707,_T_6722,_T_6721,_T_7317}; // @[Mux.scala 19:72:@4119.4]
  assign _T_7327 = _T_4267 ? _T_7325 : 16'h0; // @[Mux.scala 19:72:@4120.4]
  assign _T_7334 = {_T_6791,_T_6790,_T_6789,_T_6788,_T_6787,_T_6786,_T_6785,_T_6784}; // @[Mux.scala 19:72:@4127.4]
  assign _T_7342 = {_T_6783,_T_6782,_T_6781,_T_6780,_T_6779,_T_6794,_T_6793,_T_6792,_T_7334}; // @[Mux.scala 19:72:@4135.4]
  assign _T_7344 = _T_4268 ? _T_7342 : 16'h0; // @[Mux.scala 19:72:@4136.4]
  assign _T_7351 = {_T_6862,_T_6861,_T_6860,_T_6859,_T_6858,_T_6857,_T_6856,_T_6855}; // @[Mux.scala 19:72:@4143.4]
  assign _T_7359 = {_T_6854,_T_6853,_T_6852,_T_6851,_T_6866,_T_6865,_T_6864,_T_6863,_T_7351}; // @[Mux.scala 19:72:@4151.4]
  assign _T_7361 = _T_4269 ? _T_7359 : 16'h0; // @[Mux.scala 19:72:@4152.4]
  assign _T_7368 = {_T_6933,_T_6932,_T_6931,_T_6930,_T_6929,_T_6928,_T_6927,_T_6926}; // @[Mux.scala 19:72:@4159.4]
  assign _T_7376 = {_T_6925,_T_6924,_T_6923,_T_6938,_T_6937,_T_6936,_T_6935,_T_6934,_T_7368}; // @[Mux.scala 19:72:@4167.4]
  assign _T_7378 = _T_4270 ? _T_7376 : 16'h0; // @[Mux.scala 19:72:@4168.4]
  assign _T_7385 = {_T_7004,_T_7003,_T_7002,_T_7001,_T_7000,_T_6999,_T_6998,_T_6997}; // @[Mux.scala 19:72:@4175.4]
  assign _T_7393 = {_T_6996,_T_6995,_T_7010,_T_7009,_T_7008,_T_7007,_T_7006,_T_7005,_T_7385}; // @[Mux.scala 19:72:@4183.4]
  assign _T_7395 = _T_4271 ? _T_7393 : 16'h0; // @[Mux.scala 19:72:@4184.4]
  assign _T_7402 = {_T_7075,_T_7074,_T_7073,_T_7072,_T_7071,_T_7070,_T_7069,_T_7068}; // @[Mux.scala 19:72:@4191.4]
  assign _T_7410 = {_T_7067,_T_7082,_T_7081,_T_7080,_T_7079,_T_7078,_T_7077,_T_7076,_T_7402}; // @[Mux.scala 19:72:@4199.4]
  assign _T_7412 = _T_4272 ? _T_7410 : 16'h0; // @[Mux.scala 19:72:@4200.4]
  assign _T_7413 = _T_7157 | _T_7174; // @[Mux.scala 19:72:@4201.4]
  assign _T_7414 = _T_7413 | _T_7191; // @[Mux.scala 19:72:@4202.4]
  assign _T_7415 = _T_7414 | _T_7208; // @[Mux.scala 19:72:@4203.4]
  assign _T_7416 = _T_7415 | _T_7225; // @[Mux.scala 19:72:@4204.4]
  assign _T_7417 = _T_7416 | _T_7242; // @[Mux.scala 19:72:@4205.4]
  assign _T_7418 = _T_7417 | _T_7259; // @[Mux.scala 19:72:@4206.4]
  assign _T_7419 = _T_7418 | _T_7276; // @[Mux.scala 19:72:@4207.4]
  assign _T_7420 = _T_7419 | _T_7293; // @[Mux.scala 19:72:@4208.4]
  assign _T_7421 = _T_7420 | _T_7310; // @[Mux.scala 19:72:@4209.4]
  assign _T_7422 = _T_7421 | _T_7327; // @[Mux.scala 19:72:@4210.4]
  assign _T_7423 = _T_7422 | _T_7344; // @[Mux.scala 19:72:@4211.4]
  assign _T_7424 = _T_7423 | _T_7361; // @[Mux.scala 19:72:@4212.4]
  assign _T_7425 = _T_7424 | _T_7378; // @[Mux.scala 19:72:@4213.4]
  assign _T_7426 = _T_7425 | _T_7395; // @[Mux.scala 19:72:@4214.4]
  assign _T_7427 = _T_7426 | _T_7412; // @[Mux.scala 19:72:@4215.4]
  assign inputDataPriorityPorts_0_0 = _T_7427[0]; // @[Mux.scala 19:72:@4219.4]
  assign inputDataPriorityPorts_0_1 = _T_7427[1]; // @[Mux.scala 19:72:@4221.4]
  assign inputDataPriorityPorts_0_2 = _T_7427[2]; // @[Mux.scala 19:72:@4223.4]
  assign inputDataPriorityPorts_0_3 = _T_7427[3]; // @[Mux.scala 19:72:@4225.4]
  assign inputDataPriorityPorts_0_4 = _T_7427[4]; // @[Mux.scala 19:72:@4227.4]
  assign inputDataPriorityPorts_0_5 = _T_7427[5]; // @[Mux.scala 19:72:@4229.4]
  assign inputDataPriorityPorts_0_6 = _T_7427[6]; // @[Mux.scala 19:72:@4231.4]
  assign inputDataPriorityPorts_0_7 = _T_7427[7]; // @[Mux.scala 19:72:@4233.4]
  assign inputDataPriorityPorts_0_8 = _T_7427[8]; // @[Mux.scala 19:72:@4235.4]
  assign inputDataPriorityPorts_0_9 = _T_7427[9]; // @[Mux.scala 19:72:@4237.4]
  assign inputDataPriorityPorts_0_10 = _T_7427[10]; // @[Mux.scala 19:72:@4239.4]
  assign inputDataPriorityPorts_0_11 = _T_7427[11]; // @[Mux.scala 19:72:@4241.4]
  assign inputDataPriorityPorts_0_12 = _T_7427[12]; // @[Mux.scala 19:72:@4243.4]
  assign inputDataPriorityPorts_0_13 = _T_7427[13]; // @[Mux.scala 19:72:@4245.4]
  assign inputDataPriorityPorts_0_14 = _T_7427[14]; // @[Mux.scala 19:72:@4247.4]
  assign inputDataPriorityPorts_0_15 = _T_7427[15]; // @[Mux.scala 19:72:@4249.4]
  assign _T_7573 = inputAddrPriorityPorts_0_0 & _T_4114; // @[AxiStoreQueue.scala 214:52:@4273.6]
  assign _T_7574 = _T_7573 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4274.6]
  assign _GEN_992 = _T_7574 ? io_addressFromStorePorts_0 : addrQ_0; // @[AxiStoreQueue.scala 215:40:@4278.6]
  assign _GEN_993 = _T_7574 ? 1'h1 : addrKnown_0; // @[AxiStoreQueue.scala 215:40:@4278.6]
  assign _T_7590 = inputDataPriorityPorts_0_0 & _T_4184; // @[AxiStoreQueue.scala 220:52:@4283.6]
  assign _T_7591 = _T_7590 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4284.6]
  assign _GEN_994 = _T_7591 ? io_dataFromStorePorts_0 : dataQ_0; // @[AxiStoreQueue.scala 221:40:@4288.6]
  assign _GEN_995 = _T_7591 ? 1'h1 : dataKnown_0; // @[AxiStoreQueue.scala 221:40:@4288.6]
  assign _GEN_996 = initBits_0 ? 1'h0 : _GEN_993; // @[AxiStoreQueue.scala 209:35:@4267.4]
  assign _GEN_997 = initBits_0 ? 1'h0 : _GEN_995; // @[AxiStoreQueue.scala 209:35:@4267.4]
  assign _GEN_998 = initBits_0 ? addrQ_0 : _GEN_992; // @[AxiStoreQueue.scala 209:35:@4267.4]
  assign _GEN_999 = initBits_0 ? dataQ_0 : _GEN_994; // @[AxiStoreQueue.scala 209:35:@4267.4]
  assign _T_7609 = inputAddrPriorityPorts_0_1 & _T_4117; // @[AxiStoreQueue.scala 214:52:@4299.6]
  assign _T_7610 = _T_7609 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4300.6]
  assign _GEN_1000 = _T_7610 ? io_addressFromStorePorts_0 : addrQ_1; // @[AxiStoreQueue.scala 215:40:@4304.6]
  assign _GEN_1001 = _T_7610 ? 1'h1 : addrKnown_1; // @[AxiStoreQueue.scala 215:40:@4304.6]
  assign _T_7626 = inputDataPriorityPorts_0_1 & _T_4187; // @[AxiStoreQueue.scala 220:52:@4309.6]
  assign _T_7627 = _T_7626 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4310.6]
  assign _GEN_1002 = _T_7627 ? io_dataFromStorePorts_0 : dataQ_1; // @[AxiStoreQueue.scala 221:40:@4314.6]
  assign _GEN_1003 = _T_7627 ? 1'h1 : dataKnown_1; // @[AxiStoreQueue.scala 221:40:@4314.6]
  assign _GEN_1004 = initBits_1 ? 1'h0 : _GEN_1001; // @[AxiStoreQueue.scala 209:35:@4293.4]
  assign _GEN_1005 = initBits_1 ? 1'h0 : _GEN_1003; // @[AxiStoreQueue.scala 209:35:@4293.4]
  assign _GEN_1006 = initBits_1 ? addrQ_1 : _GEN_1000; // @[AxiStoreQueue.scala 209:35:@4293.4]
  assign _GEN_1007 = initBits_1 ? dataQ_1 : _GEN_1002; // @[AxiStoreQueue.scala 209:35:@4293.4]
  assign _T_7645 = inputAddrPriorityPorts_0_2 & _T_4120; // @[AxiStoreQueue.scala 214:52:@4325.6]
  assign _T_7646 = _T_7645 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4326.6]
  assign _GEN_1008 = _T_7646 ? io_addressFromStorePorts_0 : addrQ_2; // @[AxiStoreQueue.scala 215:40:@4330.6]
  assign _GEN_1009 = _T_7646 ? 1'h1 : addrKnown_2; // @[AxiStoreQueue.scala 215:40:@4330.6]
  assign _T_7662 = inputDataPriorityPorts_0_2 & _T_4190; // @[AxiStoreQueue.scala 220:52:@4335.6]
  assign _T_7663 = _T_7662 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4336.6]
  assign _GEN_1010 = _T_7663 ? io_dataFromStorePorts_0 : dataQ_2; // @[AxiStoreQueue.scala 221:40:@4340.6]
  assign _GEN_1011 = _T_7663 ? 1'h1 : dataKnown_2; // @[AxiStoreQueue.scala 221:40:@4340.6]
  assign _GEN_1012 = initBits_2 ? 1'h0 : _GEN_1009; // @[AxiStoreQueue.scala 209:35:@4319.4]
  assign _GEN_1013 = initBits_2 ? 1'h0 : _GEN_1011; // @[AxiStoreQueue.scala 209:35:@4319.4]
  assign _GEN_1014 = initBits_2 ? addrQ_2 : _GEN_1008; // @[AxiStoreQueue.scala 209:35:@4319.4]
  assign _GEN_1015 = initBits_2 ? dataQ_2 : _GEN_1010; // @[AxiStoreQueue.scala 209:35:@4319.4]
  assign _T_7681 = inputAddrPriorityPorts_0_3 & _T_4123; // @[AxiStoreQueue.scala 214:52:@4351.6]
  assign _T_7682 = _T_7681 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4352.6]
  assign _GEN_1016 = _T_7682 ? io_addressFromStorePorts_0 : addrQ_3; // @[AxiStoreQueue.scala 215:40:@4356.6]
  assign _GEN_1017 = _T_7682 ? 1'h1 : addrKnown_3; // @[AxiStoreQueue.scala 215:40:@4356.6]
  assign _T_7698 = inputDataPriorityPorts_0_3 & _T_4193; // @[AxiStoreQueue.scala 220:52:@4361.6]
  assign _T_7699 = _T_7698 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4362.6]
  assign _GEN_1018 = _T_7699 ? io_dataFromStorePorts_0 : dataQ_3; // @[AxiStoreQueue.scala 221:40:@4366.6]
  assign _GEN_1019 = _T_7699 ? 1'h1 : dataKnown_3; // @[AxiStoreQueue.scala 221:40:@4366.6]
  assign _GEN_1020 = initBits_3 ? 1'h0 : _GEN_1017; // @[AxiStoreQueue.scala 209:35:@4345.4]
  assign _GEN_1021 = initBits_3 ? 1'h0 : _GEN_1019; // @[AxiStoreQueue.scala 209:35:@4345.4]
  assign _GEN_1022 = initBits_3 ? addrQ_3 : _GEN_1016; // @[AxiStoreQueue.scala 209:35:@4345.4]
  assign _GEN_1023 = initBits_3 ? dataQ_3 : _GEN_1018; // @[AxiStoreQueue.scala 209:35:@4345.4]
  assign _T_7717 = inputAddrPriorityPorts_0_4 & _T_4126; // @[AxiStoreQueue.scala 214:52:@4377.6]
  assign _T_7718 = _T_7717 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4378.6]
  assign _GEN_1024 = _T_7718 ? io_addressFromStorePorts_0 : addrQ_4; // @[AxiStoreQueue.scala 215:40:@4382.6]
  assign _GEN_1025 = _T_7718 ? 1'h1 : addrKnown_4; // @[AxiStoreQueue.scala 215:40:@4382.6]
  assign _T_7734 = inputDataPriorityPorts_0_4 & _T_4196; // @[AxiStoreQueue.scala 220:52:@4387.6]
  assign _T_7735 = _T_7734 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4388.6]
  assign _GEN_1026 = _T_7735 ? io_dataFromStorePorts_0 : dataQ_4; // @[AxiStoreQueue.scala 221:40:@4392.6]
  assign _GEN_1027 = _T_7735 ? 1'h1 : dataKnown_4; // @[AxiStoreQueue.scala 221:40:@4392.6]
  assign _GEN_1028 = initBits_4 ? 1'h0 : _GEN_1025; // @[AxiStoreQueue.scala 209:35:@4371.4]
  assign _GEN_1029 = initBits_4 ? 1'h0 : _GEN_1027; // @[AxiStoreQueue.scala 209:35:@4371.4]
  assign _GEN_1030 = initBits_4 ? addrQ_4 : _GEN_1024; // @[AxiStoreQueue.scala 209:35:@4371.4]
  assign _GEN_1031 = initBits_4 ? dataQ_4 : _GEN_1026; // @[AxiStoreQueue.scala 209:35:@4371.4]
  assign _T_7753 = inputAddrPriorityPorts_0_5 & _T_4129; // @[AxiStoreQueue.scala 214:52:@4403.6]
  assign _T_7754 = _T_7753 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4404.6]
  assign _GEN_1032 = _T_7754 ? io_addressFromStorePorts_0 : addrQ_5; // @[AxiStoreQueue.scala 215:40:@4408.6]
  assign _GEN_1033 = _T_7754 ? 1'h1 : addrKnown_5; // @[AxiStoreQueue.scala 215:40:@4408.6]
  assign _T_7770 = inputDataPriorityPorts_0_5 & _T_4199; // @[AxiStoreQueue.scala 220:52:@4413.6]
  assign _T_7771 = _T_7770 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4414.6]
  assign _GEN_1034 = _T_7771 ? io_dataFromStorePorts_0 : dataQ_5; // @[AxiStoreQueue.scala 221:40:@4418.6]
  assign _GEN_1035 = _T_7771 ? 1'h1 : dataKnown_5; // @[AxiStoreQueue.scala 221:40:@4418.6]
  assign _GEN_1036 = initBits_5 ? 1'h0 : _GEN_1033; // @[AxiStoreQueue.scala 209:35:@4397.4]
  assign _GEN_1037 = initBits_5 ? 1'h0 : _GEN_1035; // @[AxiStoreQueue.scala 209:35:@4397.4]
  assign _GEN_1038 = initBits_5 ? addrQ_5 : _GEN_1032; // @[AxiStoreQueue.scala 209:35:@4397.4]
  assign _GEN_1039 = initBits_5 ? dataQ_5 : _GEN_1034; // @[AxiStoreQueue.scala 209:35:@4397.4]
  assign _T_7789 = inputAddrPriorityPorts_0_6 & _T_4132; // @[AxiStoreQueue.scala 214:52:@4429.6]
  assign _T_7790 = _T_7789 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4430.6]
  assign _GEN_1040 = _T_7790 ? io_addressFromStorePorts_0 : addrQ_6; // @[AxiStoreQueue.scala 215:40:@4434.6]
  assign _GEN_1041 = _T_7790 ? 1'h1 : addrKnown_6; // @[AxiStoreQueue.scala 215:40:@4434.6]
  assign _T_7806 = inputDataPriorityPorts_0_6 & _T_4202; // @[AxiStoreQueue.scala 220:52:@4439.6]
  assign _T_7807 = _T_7806 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4440.6]
  assign _GEN_1042 = _T_7807 ? io_dataFromStorePorts_0 : dataQ_6; // @[AxiStoreQueue.scala 221:40:@4444.6]
  assign _GEN_1043 = _T_7807 ? 1'h1 : dataKnown_6; // @[AxiStoreQueue.scala 221:40:@4444.6]
  assign _GEN_1044 = initBits_6 ? 1'h0 : _GEN_1041; // @[AxiStoreQueue.scala 209:35:@4423.4]
  assign _GEN_1045 = initBits_6 ? 1'h0 : _GEN_1043; // @[AxiStoreQueue.scala 209:35:@4423.4]
  assign _GEN_1046 = initBits_6 ? addrQ_6 : _GEN_1040; // @[AxiStoreQueue.scala 209:35:@4423.4]
  assign _GEN_1047 = initBits_6 ? dataQ_6 : _GEN_1042; // @[AxiStoreQueue.scala 209:35:@4423.4]
  assign _T_7825 = inputAddrPriorityPorts_0_7 & _T_4135; // @[AxiStoreQueue.scala 214:52:@4455.6]
  assign _T_7826 = _T_7825 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4456.6]
  assign _GEN_1048 = _T_7826 ? io_addressFromStorePorts_0 : addrQ_7; // @[AxiStoreQueue.scala 215:40:@4460.6]
  assign _GEN_1049 = _T_7826 ? 1'h1 : addrKnown_7; // @[AxiStoreQueue.scala 215:40:@4460.6]
  assign _T_7842 = inputDataPriorityPorts_0_7 & _T_4205; // @[AxiStoreQueue.scala 220:52:@4465.6]
  assign _T_7843 = _T_7842 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4466.6]
  assign _GEN_1050 = _T_7843 ? io_dataFromStorePorts_0 : dataQ_7; // @[AxiStoreQueue.scala 221:40:@4470.6]
  assign _GEN_1051 = _T_7843 ? 1'h1 : dataKnown_7; // @[AxiStoreQueue.scala 221:40:@4470.6]
  assign _GEN_1052 = initBits_7 ? 1'h0 : _GEN_1049; // @[AxiStoreQueue.scala 209:35:@4449.4]
  assign _GEN_1053 = initBits_7 ? 1'h0 : _GEN_1051; // @[AxiStoreQueue.scala 209:35:@4449.4]
  assign _GEN_1054 = initBits_7 ? addrQ_7 : _GEN_1048; // @[AxiStoreQueue.scala 209:35:@4449.4]
  assign _GEN_1055 = initBits_7 ? dataQ_7 : _GEN_1050; // @[AxiStoreQueue.scala 209:35:@4449.4]
  assign _T_7861 = inputAddrPriorityPorts_0_8 & _T_4138; // @[AxiStoreQueue.scala 214:52:@4481.6]
  assign _T_7862 = _T_7861 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4482.6]
  assign _GEN_1056 = _T_7862 ? io_addressFromStorePorts_0 : addrQ_8; // @[AxiStoreQueue.scala 215:40:@4486.6]
  assign _GEN_1057 = _T_7862 ? 1'h1 : addrKnown_8; // @[AxiStoreQueue.scala 215:40:@4486.6]
  assign _T_7878 = inputDataPriorityPorts_0_8 & _T_4208; // @[AxiStoreQueue.scala 220:52:@4491.6]
  assign _T_7879 = _T_7878 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4492.6]
  assign _GEN_1058 = _T_7879 ? io_dataFromStorePorts_0 : dataQ_8; // @[AxiStoreQueue.scala 221:40:@4496.6]
  assign _GEN_1059 = _T_7879 ? 1'h1 : dataKnown_8; // @[AxiStoreQueue.scala 221:40:@4496.6]
  assign _GEN_1060 = initBits_8 ? 1'h0 : _GEN_1057; // @[AxiStoreQueue.scala 209:35:@4475.4]
  assign _GEN_1061 = initBits_8 ? 1'h0 : _GEN_1059; // @[AxiStoreQueue.scala 209:35:@4475.4]
  assign _GEN_1062 = initBits_8 ? addrQ_8 : _GEN_1056; // @[AxiStoreQueue.scala 209:35:@4475.4]
  assign _GEN_1063 = initBits_8 ? dataQ_8 : _GEN_1058; // @[AxiStoreQueue.scala 209:35:@4475.4]
  assign _T_7897 = inputAddrPriorityPorts_0_9 & _T_4141; // @[AxiStoreQueue.scala 214:52:@4507.6]
  assign _T_7898 = _T_7897 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4508.6]
  assign _GEN_1064 = _T_7898 ? io_addressFromStorePorts_0 : addrQ_9; // @[AxiStoreQueue.scala 215:40:@4512.6]
  assign _GEN_1065 = _T_7898 ? 1'h1 : addrKnown_9; // @[AxiStoreQueue.scala 215:40:@4512.6]
  assign _T_7914 = inputDataPriorityPorts_0_9 & _T_4211; // @[AxiStoreQueue.scala 220:52:@4517.6]
  assign _T_7915 = _T_7914 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4518.6]
  assign _GEN_1066 = _T_7915 ? io_dataFromStorePorts_0 : dataQ_9; // @[AxiStoreQueue.scala 221:40:@4522.6]
  assign _GEN_1067 = _T_7915 ? 1'h1 : dataKnown_9; // @[AxiStoreQueue.scala 221:40:@4522.6]
  assign _GEN_1068 = initBits_9 ? 1'h0 : _GEN_1065; // @[AxiStoreQueue.scala 209:35:@4501.4]
  assign _GEN_1069 = initBits_9 ? 1'h0 : _GEN_1067; // @[AxiStoreQueue.scala 209:35:@4501.4]
  assign _GEN_1070 = initBits_9 ? addrQ_9 : _GEN_1064; // @[AxiStoreQueue.scala 209:35:@4501.4]
  assign _GEN_1071 = initBits_9 ? dataQ_9 : _GEN_1066; // @[AxiStoreQueue.scala 209:35:@4501.4]
  assign _T_7933 = inputAddrPriorityPorts_0_10 & _T_4144; // @[AxiStoreQueue.scala 214:52:@4533.6]
  assign _T_7934 = _T_7933 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4534.6]
  assign _GEN_1072 = _T_7934 ? io_addressFromStorePorts_0 : addrQ_10; // @[AxiStoreQueue.scala 215:40:@4538.6]
  assign _GEN_1073 = _T_7934 ? 1'h1 : addrKnown_10; // @[AxiStoreQueue.scala 215:40:@4538.6]
  assign _T_7950 = inputDataPriorityPorts_0_10 & _T_4214; // @[AxiStoreQueue.scala 220:52:@4543.6]
  assign _T_7951 = _T_7950 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4544.6]
  assign _GEN_1074 = _T_7951 ? io_dataFromStorePorts_0 : dataQ_10; // @[AxiStoreQueue.scala 221:40:@4548.6]
  assign _GEN_1075 = _T_7951 ? 1'h1 : dataKnown_10; // @[AxiStoreQueue.scala 221:40:@4548.6]
  assign _GEN_1076 = initBits_10 ? 1'h0 : _GEN_1073; // @[AxiStoreQueue.scala 209:35:@4527.4]
  assign _GEN_1077 = initBits_10 ? 1'h0 : _GEN_1075; // @[AxiStoreQueue.scala 209:35:@4527.4]
  assign _GEN_1078 = initBits_10 ? addrQ_10 : _GEN_1072; // @[AxiStoreQueue.scala 209:35:@4527.4]
  assign _GEN_1079 = initBits_10 ? dataQ_10 : _GEN_1074; // @[AxiStoreQueue.scala 209:35:@4527.4]
  assign _T_7969 = inputAddrPriorityPorts_0_11 & _T_4147; // @[AxiStoreQueue.scala 214:52:@4559.6]
  assign _T_7970 = _T_7969 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4560.6]
  assign _GEN_1080 = _T_7970 ? io_addressFromStorePorts_0 : addrQ_11; // @[AxiStoreQueue.scala 215:40:@4564.6]
  assign _GEN_1081 = _T_7970 ? 1'h1 : addrKnown_11; // @[AxiStoreQueue.scala 215:40:@4564.6]
  assign _T_7986 = inputDataPriorityPorts_0_11 & _T_4217; // @[AxiStoreQueue.scala 220:52:@4569.6]
  assign _T_7987 = _T_7986 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4570.6]
  assign _GEN_1082 = _T_7987 ? io_dataFromStorePorts_0 : dataQ_11; // @[AxiStoreQueue.scala 221:40:@4574.6]
  assign _GEN_1083 = _T_7987 ? 1'h1 : dataKnown_11; // @[AxiStoreQueue.scala 221:40:@4574.6]
  assign _GEN_1084 = initBits_11 ? 1'h0 : _GEN_1081; // @[AxiStoreQueue.scala 209:35:@4553.4]
  assign _GEN_1085 = initBits_11 ? 1'h0 : _GEN_1083; // @[AxiStoreQueue.scala 209:35:@4553.4]
  assign _GEN_1086 = initBits_11 ? addrQ_11 : _GEN_1080; // @[AxiStoreQueue.scala 209:35:@4553.4]
  assign _GEN_1087 = initBits_11 ? dataQ_11 : _GEN_1082; // @[AxiStoreQueue.scala 209:35:@4553.4]
  assign _T_8005 = inputAddrPriorityPorts_0_12 & _T_4150; // @[AxiStoreQueue.scala 214:52:@4585.6]
  assign _T_8006 = _T_8005 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4586.6]
  assign _GEN_1088 = _T_8006 ? io_addressFromStorePorts_0 : addrQ_12; // @[AxiStoreQueue.scala 215:40:@4590.6]
  assign _GEN_1089 = _T_8006 ? 1'h1 : addrKnown_12; // @[AxiStoreQueue.scala 215:40:@4590.6]
  assign _T_8022 = inputDataPriorityPorts_0_12 & _T_4220; // @[AxiStoreQueue.scala 220:52:@4595.6]
  assign _T_8023 = _T_8022 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4596.6]
  assign _GEN_1090 = _T_8023 ? io_dataFromStorePorts_0 : dataQ_12; // @[AxiStoreQueue.scala 221:40:@4600.6]
  assign _GEN_1091 = _T_8023 ? 1'h1 : dataKnown_12; // @[AxiStoreQueue.scala 221:40:@4600.6]
  assign _GEN_1092 = initBits_12 ? 1'h0 : _GEN_1089; // @[AxiStoreQueue.scala 209:35:@4579.4]
  assign _GEN_1093 = initBits_12 ? 1'h0 : _GEN_1091; // @[AxiStoreQueue.scala 209:35:@4579.4]
  assign _GEN_1094 = initBits_12 ? addrQ_12 : _GEN_1088; // @[AxiStoreQueue.scala 209:35:@4579.4]
  assign _GEN_1095 = initBits_12 ? dataQ_12 : _GEN_1090; // @[AxiStoreQueue.scala 209:35:@4579.4]
  assign _T_8041 = inputAddrPriorityPorts_0_13 & _T_4153; // @[AxiStoreQueue.scala 214:52:@4611.6]
  assign _T_8042 = _T_8041 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4612.6]
  assign _GEN_1096 = _T_8042 ? io_addressFromStorePorts_0 : addrQ_13; // @[AxiStoreQueue.scala 215:40:@4616.6]
  assign _GEN_1097 = _T_8042 ? 1'h1 : addrKnown_13; // @[AxiStoreQueue.scala 215:40:@4616.6]
  assign _T_8058 = inputDataPriorityPorts_0_13 & _T_4223; // @[AxiStoreQueue.scala 220:52:@4621.6]
  assign _T_8059 = _T_8058 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4622.6]
  assign _GEN_1098 = _T_8059 ? io_dataFromStorePorts_0 : dataQ_13; // @[AxiStoreQueue.scala 221:40:@4626.6]
  assign _GEN_1099 = _T_8059 ? 1'h1 : dataKnown_13; // @[AxiStoreQueue.scala 221:40:@4626.6]
  assign _GEN_1100 = initBits_13 ? 1'h0 : _GEN_1097; // @[AxiStoreQueue.scala 209:35:@4605.4]
  assign _GEN_1101 = initBits_13 ? 1'h0 : _GEN_1099; // @[AxiStoreQueue.scala 209:35:@4605.4]
  assign _GEN_1102 = initBits_13 ? addrQ_13 : _GEN_1096; // @[AxiStoreQueue.scala 209:35:@4605.4]
  assign _GEN_1103 = initBits_13 ? dataQ_13 : _GEN_1098; // @[AxiStoreQueue.scala 209:35:@4605.4]
  assign _T_8077 = inputAddrPriorityPorts_0_14 & _T_4156; // @[AxiStoreQueue.scala 214:52:@4637.6]
  assign _T_8078 = _T_8077 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4638.6]
  assign _GEN_1104 = _T_8078 ? io_addressFromStorePorts_0 : addrQ_14; // @[AxiStoreQueue.scala 215:40:@4642.6]
  assign _GEN_1105 = _T_8078 ? 1'h1 : addrKnown_14; // @[AxiStoreQueue.scala 215:40:@4642.6]
  assign _T_8094 = inputDataPriorityPorts_0_14 & _T_4226; // @[AxiStoreQueue.scala 220:52:@4647.6]
  assign _T_8095 = _T_8094 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4648.6]
  assign _GEN_1106 = _T_8095 ? io_dataFromStorePorts_0 : dataQ_14; // @[AxiStoreQueue.scala 221:40:@4652.6]
  assign _GEN_1107 = _T_8095 ? 1'h1 : dataKnown_14; // @[AxiStoreQueue.scala 221:40:@4652.6]
  assign _GEN_1108 = initBits_14 ? 1'h0 : _GEN_1105; // @[AxiStoreQueue.scala 209:35:@4631.4]
  assign _GEN_1109 = initBits_14 ? 1'h0 : _GEN_1107; // @[AxiStoreQueue.scala 209:35:@4631.4]
  assign _GEN_1110 = initBits_14 ? addrQ_14 : _GEN_1104; // @[AxiStoreQueue.scala 209:35:@4631.4]
  assign _GEN_1111 = initBits_14 ? dataQ_14 : _GEN_1106; // @[AxiStoreQueue.scala 209:35:@4631.4]
  assign _T_8113 = inputAddrPriorityPorts_0_15 & _T_4159; // @[AxiStoreQueue.scala 214:52:@4663.6]
  assign _T_8114 = _T_8113 & io_storeAddrEnable_0; // @[AxiStoreQueue.scala 214:81:@4664.6]
  assign _GEN_1112 = _T_8114 ? io_addressFromStorePorts_0 : addrQ_15; // @[AxiStoreQueue.scala 215:40:@4668.6]
  assign _GEN_1113 = _T_8114 ? 1'h1 : addrKnown_15; // @[AxiStoreQueue.scala 215:40:@4668.6]
  assign _T_8130 = inputDataPriorityPorts_0_15 & _T_4229; // @[AxiStoreQueue.scala 220:52:@4673.6]
  assign _T_8131 = _T_8130 & io_storeDataEnable_0; // @[AxiStoreQueue.scala 220:81:@4674.6]
  assign _GEN_1114 = _T_8131 ? io_dataFromStorePorts_0 : dataQ_15; // @[AxiStoreQueue.scala 221:40:@4678.6]
  assign _GEN_1115 = _T_8131 ? 1'h1 : dataKnown_15; // @[AxiStoreQueue.scala 221:40:@4678.6]
  assign _GEN_1116 = initBits_15 ? 1'h0 : _GEN_1113; // @[AxiStoreQueue.scala 209:35:@4657.4]
  assign _GEN_1117 = initBits_15 ? 1'h0 : _GEN_1115; // @[AxiStoreQueue.scala 209:35:@4657.4]
  assign _GEN_1118 = initBits_15 ? addrQ_15 : _GEN_1112; // @[AxiStoreQueue.scala 209:35:@4657.4]
  assign _GEN_1119 = initBits_15 ? dataQ_15 : _GEN_1114; // @[AxiStoreQueue.scala 209:35:@4657.4]
  assign _T_8145 = io_storeQIdxOut_ready & storeRequest; // @[AxiStoreQueue.scala 234:30:@4683.4]
  assign _T_8148 = dummyHead + 4'h1; // @[util.scala 10:8:@4685.6]
  assign _GEN_64 = _T_8148 % 5'h10; // @[util.scala 10:14:@4686.6]
  assign _T_8149 = _GEN_64[4:0]; // @[util.scala 10:14:@4686.6]
  assign _GEN_1120 = _T_8145 ? _T_8149 : {{1'd0}, dummyHead}; // @[AxiStoreQueue.scala 234:47:@4684.4]
  assign _GEN_1251 = {{3'd0}, io_bbNumStores}; // @[util.scala 10:8:@4698.6]
  assign _T_8161 = tail + _GEN_1251; // @[util.scala 10:8:@4698.6]
  assign _GEN_65 = _T_8161 % 5'h10; // @[util.scala 10:14:@4699.6]
  assign _T_8162 = _GEN_65[4:0]; // @[util.scala 10:14:@4699.6]
  assign _GEN_1138 = io_bbStart ? _T_8162 : {{1'd0}, tail}; // @[AxiStoreQueue.scala 243:20:@4697.4]
  assign _T_8164 = allocatedEntries_0 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4702.4]
  assign _T_8165 = storeCompleted_0 | _T_8164; // @[AxiStoreQueue.scala 247:81:@4703.4]
  assign _T_8167 = allocatedEntries_1 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4704.4]
  assign _T_8168 = storeCompleted_1 | _T_8167; // @[AxiStoreQueue.scala 247:81:@4705.4]
  assign _T_8170 = allocatedEntries_2 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4706.4]
  assign _T_8171 = storeCompleted_2 | _T_8170; // @[AxiStoreQueue.scala 247:81:@4707.4]
  assign _T_8173 = allocatedEntries_3 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4708.4]
  assign _T_8174 = storeCompleted_3 | _T_8173; // @[AxiStoreQueue.scala 247:81:@4709.4]
  assign _T_8176 = allocatedEntries_4 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4710.4]
  assign _T_8177 = storeCompleted_4 | _T_8176; // @[AxiStoreQueue.scala 247:81:@4711.4]
  assign _T_8179 = allocatedEntries_5 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4712.4]
  assign _T_8180 = storeCompleted_5 | _T_8179; // @[AxiStoreQueue.scala 247:81:@4713.4]
  assign _T_8182 = allocatedEntries_6 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4714.4]
  assign _T_8183 = storeCompleted_6 | _T_8182; // @[AxiStoreQueue.scala 247:81:@4715.4]
  assign _T_8185 = allocatedEntries_7 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4716.4]
  assign _T_8186 = storeCompleted_7 | _T_8185; // @[AxiStoreQueue.scala 247:81:@4717.4]
  assign _T_8188 = allocatedEntries_8 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4718.4]
  assign _T_8189 = storeCompleted_8 | _T_8188; // @[AxiStoreQueue.scala 247:81:@4719.4]
  assign _T_8191 = allocatedEntries_9 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4720.4]
  assign _T_8192 = storeCompleted_9 | _T_8191; // @[AxiStoreQueue.scala 247:81:@4721.4]
  assign _T_8194 = allocatedEntries_10 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4722.4]
  assign _T_8195 = storeCompleted_10 | _T_8194; // @[AxiStoreQueue.scala 247:81:@4723.4]
  assign _T_8197 = allocatedEntries_11 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4724.4]
  assign _T_8198 = storeCompleted_11 | _T_8197; // @[AxiStoreQueue.scala 247:81:@4725.4]
  assign _T_8200 = allocatedEntries_12 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4726.4]
  assign _T_8201 = storeCompleted_12 | _T_8200; // @[AxiStoreQueue.scala 247:81:@4727.4]
  assign _T_8203 = allocatedEntries_13 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4728.4]
  assign _T_8204 = storeCompleted_13 | _T_8203; // @[AxiStoreQueue.scala 247:81:@4729.4]
  assign _T_8206 = allocatedEntries_14 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4730.4]
  assign _T_8207 = storeCompleted_14 | _T_8206; // @[AxiStoreQueue.scala 247:81:@4731.4]
  assign _T_8209 = allocatedEntries_15 == 1'h0; // @[AxiStoreQueue.scala 247:84:@4732.4]
  assign _T_8210 = storeCompleted_15 | _T_8209; // @[AxiStoreQueue.scala 247:81:@4733.4]
  assign _T_8235 = _T_8165 & _T_8168; // @[AxiStoreQueue.scala 247:98:@4752.4]
  assign _T_8236 = _T_8235 & _T_8171; // @[AxiStoreQueue.scala 247:98:@4753.4]
  assign _T_8237 = _T_8236 & _T_8174; // @[AxiStoreQueue.scala 247:98:@4754.4]
  assign _T_8238 = _T_8237 & _T_8177; // @[AxiStoreQueue.scala 247:98:@4755.4]
  assign _T_8239 = _T_8238 & _T_8180; // @[AxiStoreQueue.scala 247:98:@4756.4]
  assign _T_8240 = _T_8239 & _T_8183; // @[AxiStoreQueue.scala 247:98:@4757.4]
  assign _T_8241 = _T_8240 & _T_8186; // @[AxiStoreQueue.scala 247:98:@4758.4]
  assign _T_8242 = _T_8241 & _T_8189; // @[AxiStoreQueue.scala 247:98:@4759.4]
  assign _T_8243 = _T_8242 & _T_8192; // @[AxiStoreQueue.scala 247:98:@4760.4]
  assign _T_8244 = _T_8243 & _T_8195; // @[AxiStoreQueue.scala 247:98:@4761.4]
  assign _T_8245 = _T_8244 & _T_8198; // @[AxiStoreQueue.scala 247:98:@4762.4]
  assign _T_8246 = _T_8245 & _T_8201; // @[AxiStoreQueue.scala 247:98:@4763.4]
  assign _T_8247 = _T_8246 & _T_8204; // @[AxiStoreQueue.scala 247:98:@4764.4]
  assign _T_8248 = _T_8247 & _T_8207; // @[AxiStoreQueue.scala 247:98:@4765.4]
  assign _GEN_1140 = 4'h1 == dummyHead ? dataQ_1 : dataQ_0; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1141 = 4'h2 == dummyHead ? dataQ_2 : _GEN_1140; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1142 = 4'h3 == dummyHead ? dataQ_3 : _GEN_1141; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1143 = 4'h4 == dummyHead ? dataQ_4 : _GEN_1142; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1144 = 4'h5 == dummyHead ? dataQ_5 : _GEN_1143; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1145 = 4'h6 == dummyHead ? dataQ_6 : _GEN_1144; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1146 = 4'h7 == dummyHead ? dataQ_7 : _GEN_1145; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1147 = 4'h8 == dummyHead ? dataQ_8 : _GEN_1146; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1148 = 4'h9 == dummyHead ? dataQ_9 : _GEN_1147; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1149 = 4'ha == dummyHead ? dataQ_10 : _GEN_1148; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1150 = 4'hb == dummyHead ? dataQ_11 : _GEN_1149; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1151 = 4'hc == dummyHead ? dataQ_12 : _GEN_1150; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1152 = 4'hd == dummyHead ? dataQ_13 : _GEN_1151; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign _GEN_1153 = 4'he == dummyHead ? dataQ_14 : _GEN_1152; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign io_storeTail = tail; // @[AxiStoreQueue.scala 256:16:@4769.4]
  assign io_storeHead = dummyHead; // @[AxiStoreQueue.scala 255:16:@4768.4]
  assign io_storeEmpty = _T_8248 & _T_8210; // @[AxiStoreQueue.scala 247:17:@4767.4]
  assign io_storeAddrDone_0 = addrKnown_0; // @[AxiStoreQueue.scala 260:20:@4818.4]
  assign io_storeAddrDone_1 = addrKnown_1; // @[AxiStoreQueue.scala 260:20:@4819.4]
  assign io_storeAddrDone_2 = addrKnown_2; // @[AxiStoreQueue.scala 260:20:@4820.4]
  assign io_storeAddrDone_3 = addrKnown_3; // @[AxiStoreQueue.scala 260:20:@4821.4]
  assign io_storeAddrDone_4 = addrKnown_4; // @[AxiStoreQueue.scala 260:20:@4822.4]
  assign io_storeAddrDone_5 = addrKnown_5; // @[AxiStoreQueue.scala 260:20:@4823.4]
  assign io_storeAddrDone_6 = addrKnown_6; // @[AxiStoreQueue.scala 260:20:@4824.4]
  assign io_storeAddrDone_7 = addrKnown_7; // @[AxiStoreQueue.scala 260:20:@4825.4]
  assign io_storeAddrDone_8 = addrKnown_8; // @[AxiStoreQueue.scala 260:20:@4826.4]
  assign io_storeAddrDone_9 = addrKnown_9; // @[AxiStoreQueue.scala 260:20:@4827.4]
  assign io_storeAddrDone_10 = addrKnown_10; // @[AxiStoreQueue.scala 260:20:@4828.4]
  assign io_storeAddrDone_11 = addrKnown_11; // @[AxiStoreQueue.scala 260:20:@4829.4]
  assign io_storeAddrDone_12 = addrKnown_12; // @[AxiStoreQueue.scala 260:20:@4830.4]
  assign io_storeAddrDone_13 = addrKnown_13; // @[AxiStoreQueue.scala 260:20:@4831.4]
  assign io_storeAddrDone_14 = addrKnown_14; // @[AxiStoreQueue.scala 260:20:@4832.4]
  assign io_storeAddrDone_15 = addrKnown_15; // @[AxiStoreQueue.scala 260:20:@4833.4]
  assign io_storeDataDone_0 = dataKnown_0; // @[AxiStoreQueue.scala 259:20:@4802.4]
  assign io_storeDataDone_1 = dataKnown_1; // @[AxiStoreQueue.scala 259:20:@4803.4]
  assign io_storeDataDone_2 = dataKnown_2; // @[AxiStoreQueue.scala 259:20:@4804.4]
  assign io_storeDataDone_3 = dataKnown_3; // @[AxiStoreQueue.scala 259:20:@4805.4]
  assign io_storeDataDone_4 = dataKnown_4; // @[AxiStoreQueue.scala 259:20:@4806.4]
  assign io_storeDataDone_5 = dataKnown_5; // @[AxiStoreQueue.scala 259:20:@4807.4]
  assign io_storeDataDone_6 = dataKnown_6; // @[AxiStoreQueue.scala 259:20:@4808.4]
  assign io_storeDataDone_7 = dataKnown_7; // @[AxiStoreQueue.scala 259:20:@4809.4]
  assign io_storeDataDone_8 = dataKnown_8; // @[AxiStoreQueue.scala 259:20:@4810.4]
  assign io_storeDataDone_9 = dataKnown_9; // @[AxiStoreQueue.scala 259:20:@4811.4]
  assign io_storeDataDone_10 = dataKnown_10; // @[AxiStoreQueue.scala 259:20:@4812.4]
  assign io_storeDataDone_11 = dataKnown_11; // @[AxiStoreQueue.scala 259:20:@4813.4]
  assign io_storeDataDone_12 = dataKnown_12; // @[AxiStoreQueue.scala 259:20:@4814.4]
  assign io_storeDataDone_13 = dataKnown_13; // @[AxiStoreQueue.scala 259:20:@4815.4]
  assign io_storeDataDone_14 = dataKnown_14; // @[AxiStoreQueue.scala 259:20:@4816.4]
  assign io_storeDataDone_15 = dataKnown_15; // @[AxiStoreQueue.scala 259:20:@4817.4]
  assign io_storeAddrQueue_0 = addrQ_0; // @[AxiStoreQueue.scala 257:21:@4770.4]
  assign io_storeAddrQueue_1 = addrQ_1; // @[AxiStoreQueue.scala 257:21:@4771.4]
  assign io_storeAddrQueue_2 = addrQ_2; // @[AxiStoreQueue.scala 257:21:@4772.4]
  assign io_storeAddrQueue_3 = addrQ_3; // @[AxiStoreQueue.scala 257:21:@4773.4]
  assign io_storeAddrQueue_4 = addrQ_4; // @[AxiStoreQueue.scala 257:21:@4774.4]
  assign io_storeAddrQueue_5 = addrQ_5; // @[AxiStoreQueue.scala 257:21:@4775.4]
  assign io_storeAddrQueue_6 = addrQ_6; // @[AxiStoreQueue.scala 257:21:@4776.4]
  assign io_storeAddrQueue_7 = addrQ_7; // @[AxiStoreQueue.scala 257:21:@4777.4]
  assign io_storeAddrQueue_8 = addrQ_8; // @[AxiStoreQueue.scala 257:21:@4778.4]
  assign io_storeAddrQueue_9 = addrQ_9; // @[AxiStoreQueue.scala 257:21:@4779.4]
  assign io_storeAddrQueue_10 = addrQ_10; // @[AxiStoreQueue.scala 257:21:@4780.4]
  assign io_storeAddrQueue_11 = addrQ_11; // @[AxiStoreQueue.scala 257:21:@4781.4]
  assign io_storeAddrQueue_12 = addrQ_12; // @[AxiStoreQueue.scala 257:21:@4782.4]
  assign io_storeAddrQueue_13 = addrQ_13; // @[AxiStoreQueue.scala 257:21:@4783.4]
  assign io_storeAddrQueue_14 = addrQ_14; // @[AxiStoreQueue.scala 257:21:@4784.4]
  assign io_storeAddrQueue_15 = addrQ_15; // @[AxiStoreQueue.scala 257:21:@4785.4]
  assign io_storeDataQueue_0 = dataQ_0; // @[AxiStoreQueue.scala 258:21:@4786.4]
  assign io_storeDataQueue_1 = dataQ_1; // @[AxiStoreQueue.scala 258:21:@4787.4]
  assign io_storeDataQueue_2 = dataQ_2; // @[AxiStoreQueue.scala 258:21:@4788.4]
  assign io_storeDataQueue_3 = dataQ_3; // @[AxiStoreQueue.scala 258:21:@4789.4]
  assign io_storeDataQueue_4 = dataQ_4; // @[AxiStoreQueue.scala 258:21:@4790.4]
  assign io_storeDataQueue_5 = dataQ_5; // @[AxiStoreQueue.scala 258:21:@4791.4]
  assign io_storeDataQueue_6 = dataQ_6; // @[AxiStoreQueue.scala 258:21:@4792.4]
  assign io_storeDataQueue_7 = dataQ_7; // @[AxiStoreQueue.scala 258:21:@4793.4]
  assign io_storeDataQueue_8 = dataQ_8; // @[AxiStoreQueue.scala 258:21:@4794.4]
  assign io_storeDataQueue_9 = dataQ_9; // @[AxiStoreQueue.scala 258:21:@4795.4]
  assign io_storeDataQueue_10 = dataQ_10; // @[AxiStoreQueue.scala 258:21:@4796.4]
  assign io_storeDataQueue_11 = dataQ_11; // @[AxiStoreQueue.scala 258:21:@4797.4]
  assign io_storeDataQueue_12 = dataQ_12; // @[AxiStoreQueue.scala 258:21:@4798.4]
  assign io_storeDataQueue_13 = dataQ_13; // @[AxiStoreQueue.scala 258:21:@4799.4]
  assign io_storeDataQueue_14 = dataQ_14; // @[AxiStoreQueue.scala 258:21:@4800.4]
  assign io_storeDataQueue_15 = dataQ_15; // @[AxiStoreQueue.scala 258:21:@4801.4]
  assign io_storeAddrToMem = 4'hf == dummyHead ? addrQ_15 : _GEN_910; // @[AxiStoreQueue.scala 263:21:@4836.4]
  assign io_storeDataToMem = 4'hf == dummyHead ? dataQ_15 : _GEN_1153; // @[AxiStoreQueue.scala 262:21:@4835.4]
  assign io_storeQIdxOut_valid = _T_3533 & _T_3550; // @[AxiStoreQueue.scala 261:25:@4834.4]
  assign io_storeQIdxOut_bits = dummyHead; // @[AxiStoreQueue.scala 157:24:@1705.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dummyHead = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  storeCompleted_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  storeCompleted_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  storeCompleted_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  storeCompleted_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  storeCompleted_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  storeCompleted_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  storeCompleted_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  storeCompleted_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  storeCompleted_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  storeCompleted_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  storeCompleted_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  storeCompleted_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  storeCompleted_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  storeCompleted_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  storeCompleted_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  storeCompleted_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  checkBits_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  checkBits_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  checkBits_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  checkBits_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  checkBits_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  checkBits_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  checkBits_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  checkBits_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  checkBits_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  checkBits_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  checkBits_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  checkBits_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  checkBits_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  checkBits_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  checkBits_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  checkBits_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  previousLoadHead = _RAND_146[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      dummyHead <= 4'h0;
    end else begin
      dummyHead <= _GEN_1120[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_1138[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1812) begin
          offsetQ_0 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1812) begin
            offsetQ_0 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1812) begin
              offsetQ_0 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1812) begin
                offsetQ_0 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1812) begin
                  offsetQ_0 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1812) begin
                    offsetQ_0 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1812) begin
                      offsetQ_0 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1812) begin
                        offsetQ_0 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1812) begin
                          offsetQ_0 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1812) begin
                            offsetQ_0 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1812) begin
                              offsetQ_0 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1812) begin
                                offsetQ_0 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1812) begin
                                  offsetQ_0 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1812) begin
                                    offsetQ_0 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1812) begin
                                      offsetQ_0 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1830) begin
          offsetQ_1 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1830) begin
            offsetQ_1 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1830) begin
              offsetQ_1 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1830) begin
                offsetQ_1 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1830) begin
                  offsetQ_1 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1830) begin
                    offsetQ_1 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1830) begin
                      offsetQ_1 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1830) begin
                        offsetQ_1 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1830) begin
                          offsetQ_1 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1830) begin
                            offsetQ_1 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1830) begin
                              offsetQ_1 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1830) begin
                                offsetQ_1 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1830) begin
                                  offsetQ_1 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1830) begin
                                    offsetQ_1 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1830) begin
                                      offsetQ_1 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1848) begin
          offsetQ_2 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1848) begin
            offsetQ_2 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1848) begin
              offsetQ_2 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1848) begin
                offsetQ_2 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1848) begin
                  offsetQ_2 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1848) begin
                    offsetQ_2 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1848) begin
                      offsetQ_2 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1848) begin
                        offsetQ_2 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1848) begin
                          offsetQ_2 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1848) begin
                            offsetQ_2 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1848) begin
                              offsetQ_2 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1848) begin
                                offsetQ_2 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1848) begin
                                  offsetQ_2 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1848) begin
                                    offsetQ_2 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1848) begin
                                      offsetQ_2 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1866) begin
          offsetQ_3 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1866) begin
            offsetQ_3 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1866) begin
              offsetQ_3 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1866) begin
                offsetQ_3 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1866) begin
                  offsetQ_3 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1866) begin
                    offsetQ_3 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1866) begin
                      offsetQ_3 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1866) begin
                        offsetQ_3 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1866) begin
                          offsetQ_3 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1866) begin
                            offsetQ_3 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1866) begin
                              offsetQ_3 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1866) begin
                                offsetQ_3 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1866) begin
                                  offsetQ_3 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1866) begin
                                    offsetQ_3 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1866) begin
                                      offsetQ_3 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_1884) begin
          offsetQ_4 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1884) begin
            offsetQ_4 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1884) begin
              offsetQ_4 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1884) begin
                offsetQ_4 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1884) begin
                  offsetQ_4 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1884) begin
                    offsetQ_4 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1884) begin
                      offsetQ_4 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1884) begin
                        offsetQ_4 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1884) begin
                          offsetQ_4 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1884) begin
                            offsetQ_4 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1884) begin
                              offsetQ_4 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1884) begin
                                offsetQ_4 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1884) begin
                                  offsetQ_4 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1884) begin
                                    offsetQ_4 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1884) begin
                                      offsetQ_4 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_1902) begin
          offsetQ_5 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1902) begin
            offsetQ_5 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1902) begin
              offsetQ_5 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1902) begin
                offsetQ_5 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1902) begin
                  offsetQ_5 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1902) begin
                    offsetQ_5 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1902) begin
                      offsetQ_5 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1902) begin
                        offsetQ_5 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1902) begin
                          offsetQ_5 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1902) begin
                            offsetQ_5 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1902) begin
                              offsetQ_5 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1902) begin
                                offsetQ_5 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1902) begin
                                  offsetQ_5 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1902) begin
                                    offsetQ_5 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1902) begin
                                      offsetQ_5 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_1920) begin
          offsetQ_6 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1920) begin
            offsetQ_6 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1920) begin
              offsetQ_6 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1920) begin
                offsetQ_6 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1920) begin
                  offsetQ_6 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1920) begin
                    offsetQ_6 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1920) begin
                      offsetQ_6 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1920) begin
                        offsetQ_6 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1920) begin
                          offsetQ_6 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1920) begin
                            offsetQ_6 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1920) begin
                              offsetQ_6 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1920) begin
                                offsetQ_6 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1920) begin
                                  offsetQ_6 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1920) begin
                                    offsetQ_6 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1920) begin
                                      offsetQ_6 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_1938) begin
          offsetQ_7 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1938) begin
            offsetQ_7 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1938) begin
              offsetQ_7 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1938) begin
                offsetQ_7 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1938) begin
                  offsetQ_7 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1938) begin
                    offsetQ_7 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1938) begin
                      offsetQ_7 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1938) begin
                        offsetQ_7 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1938) begin
                          offsetQ_7 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1938) begin
                            offsetQ_7 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1938) begin
                              offsetQ_7 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1938) begin
                                offsetQ_7 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1938) begin
                                  offsetQ_7 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1938) begin
                                    offsetQ_7 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1938) begin
                                      offsetQ_7 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_1956) begin
          offsetQ_8 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1956) begin
            offsetQ_8 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1956) begin
              offsetQ_8 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1956) begin
                offsetQ_8 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1956) begin
                  offsetQ_8 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1956) begin
                    offsetQ_8 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1956) begin
                      offsetQ_8 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1956) begin
                        offsetQ_8 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1956) begin
                          offsetQ_8 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1956) begin
                            offsetQ_8 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1956) begin
                              offsetQ_8 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1956) begin
                                offsetQ_8 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1956) begin
                                  offsetQ_8 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1956) begin
                                    offsetQ_8 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1956) begin
                                      offsetQ_8 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_1974) begin
          offsetQ_9 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1974) begin
            offsetQ_9 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1974) begin
              offsetQ_9 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1974) begin
                offsetQ_9 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1974) begin
                  offsetQ_9 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1974) begin
                    offsetQ_9 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1974) begin
                      offsetQ_9 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1974) begin
                        offsetQ_9 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1974) begin
                          offsetQ_9 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1974) begin
                            offsetQ_9 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1974) begin
                              offsetQ_9 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1974) begin
                                offsetQ_9 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1974) begin
                                  offsetQ_9 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1974) begin
                                    offsetQ_9 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1974) begin
                                      offsetQ_9 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_1992) begin
          offsetQ_10 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_1992) begin
            offsetQ_10 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_1992) begin
              offsetQ_10 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_1992) begin
                offsetQ_10 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_1992) begin
                  offsetQ_10 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_1992) begin
                    offsetQ_10 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_1992) begin
                      offsetQ_10 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_1992) begin
                        offsetQ_10 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_1992) begin
                          offsetQ_10 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_1992) begin
                            offsetQ_10 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_1992) begin
                              offsetQ_10 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_1992) begin
                                offsetQ_10 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_1992) begin
                                  offsetQ_10 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1992) begin
                                    offsetQ_10 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1992) begin
                                      offsetQ_10 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2010) begin
          offsetQ_11 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2010) begin
            offsetQ_11 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2010) begin
              offsetQ_11 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2010) begin
                offsetQ_11 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2010) begin
                  offsetQ_11 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2010) begin
                    offsetQ_11 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2010) begin
                      offsetQ_11 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2010) begin
                        offsetQ_11 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2010) begin
                          offsetQ_11 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2010) begin
                            offsetQ_11 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2010) begin
                              offsetQ_11 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2010) begin
                                offsetQ_11 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2010) begin
                                  offsetQ_11 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2010) begin
                                    offsetQ_11 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2010) begin
                                      offsetQ_11 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2028) begin
          offsetQ_12 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2028) begin
            offsetQ_12 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2028) begin
              offsetQ_12 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2028) begin
                offsetQ_12 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2028) begin
                  offsetQ_12 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2028) begin
                    offsetQ_12 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2028) begin
                      offsetQ_12 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2028) begin
                        offsetQ_12 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2028) begin
                          offsetQ_12 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2028) begin
                            offsetQ_12 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2028) begin
                              offsetQ_12 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2028) begin
                                offsetQ_12 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2028) begin
                                  offsetQ_12 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2028) begin
                                    offsetQ_12 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2028) begin
                                      offsetQ_12 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2046) begin
          offsetQ_13 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2046) begin
            offsetQ_13 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2046) begin
              offsetQ_13 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2046) begin
                offsetQ_13 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2046) begin
                  offsetQ_13 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2046) begin
                    offsetQ_13 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2046) begin
                      offsetQ_13 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2046) begin
                        offsetQ_13 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2046) begin
                          offsetQ_13 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2046) begin
                            offsetQ_13 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2046) begin
                              offsetQ_13 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2046) begin
                                offsetQ_13 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2046) begin
                                  offsetQ_13 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2046) begin
                                    offsetQ_13 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2046) begin
                                      offsetQ_13 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2064) begin
          offsetQ_14 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2064) begin
            offsetQ_14 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2064) begin
              offsetQ_14 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2064) begin
                offsetQ_14 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2064) begin
                  offsetQ_14 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2064) begin
                    offsetQ_14 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2064) begin
                      offsetQ_14 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2064) begin
                        offsetQ_14 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2064) begin
                          offsetQ_14 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2064) begin
                            offsetQ_14 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2064) begin
                              offsetQ_14 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2064) begin
                                offsetQ_14 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2064) begin
                                  offsetQ_14 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2064) begin
                                    offsetQ_14 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2064) begin
                                      offsetQ_14 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2082) begin
          offsetQ_15 <= io_bbStoreOffsets_15;
        end else begin
          if (4'he == _T_2082) begin
            offsetQ_15 <= io_bbStoreOffsets_14;
          end else begin
            if (4'hd == _T_2082) begin
              offsetQ_15 <= io_bbStoreOffsets_13;
            end else begin
              if (4'hc == _T_2082) begin
                offsetQ_15 <= io_bbStoreOffsets_12;
              end else begin
                if (4'hb == _T_2082) begin
                  offsetQ_15 <= io_bbStoreOffsets_11;
                end else begin
                  if (4'ha == _T_2082) begin
                    offsetQ_15 <= io_bbStoreOffsets_10;
                  end else begin
                    if (4'h9 == _T_2082) begin
                      offsetQ_15 <= io_bbStoreOffsets_9;
                    end else begin
                      if (4'h8 == _T_2082) begin
                        offsetQ_15 <= io_bbStoreOffsets_8;
                      end else begin
                        if (4'h7 == _T_2082) begin
                          offsetQ_15 <= io_bbStoreOffsets_7;
                        end else begin
                          if (4'h6 == _T_2082) begin
                            offsetQ_15 <= io_bbStoreOffsets_6;
                          end else begin
                            if (4'h5 == _T_2082) begin
                              offsetQ_15 <= io_bbStoreOffsets_5;
                            end else begin
                              if (4'h4 == _T_2082) begin
                                offsetQ_15 <= io_bbStoreOffsets_4;
                              end else begin
                                if (4'h3 == _T_2082) begin
                                  offsetQ_15 <= io_bbStoreOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2082) begin
                                    offsetQ_15 <= io_bbStoreOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2082) begin
                                      offsetQ_15 <= io_bbStoreOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbStoreOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        portQ_0 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        portQ_1 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        portQ_2 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        portQ_3 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        portQ_4 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        portQ_5 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        portQ_6 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        portQ_7 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        portQ_8 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        portQ_9 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        portQ_10 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        portQ_11 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        portQ_12 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        portQ_13 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        portQ_14 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        portQ_15 <= 1'h0;
      end
    end
    if (reset) begin
      addrQ_0 <= 31'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_7574) begin
          addrQ_0 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 31'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_7610) begin
          addrQ_1 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 31'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_7646) begin
          addrQ_2 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 31'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_7682) begin
          addrQ_3 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 31'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_7718) begin
          addrQ_4 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 31'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_7754) begin
          addrQ_5 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 31'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_7790) begin
          addrQ_6 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 31'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_7826) begin
          addrQ_7 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 31'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_7862) begin
          addrQ_8 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 31'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_7898) begin
          addrQ_9 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 31'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_7934) begin
          addrQ_10 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 31'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_7970) begin
          addrQ_11 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 31'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_8006) begin
          addrQ_12 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 31'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_8042) begin
          addrQ_13 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 31'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_8078) begin
          addrQ_14 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 31'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_8114) begin
          addrQ_15 <= io_addressFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_7591) begin
          dataQ_0 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_7627) begin
          dataQ_1 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_7663) begin
          dataQ_2 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_7699) begin
          dataQ_3 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_7735) begin
          dataQ_4 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_7771) begin
          dataQ_5 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_7807) begin
          dataQ_6 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_7843) begin
          dataQ_7 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_7879) begin
          dataQ_8 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_7915) begin
          dataQ_9 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_7951) begin
          dataQ_10 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_7987) begin
          dataQ_11 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_8023) begin
          dataQ_12 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_8059) begin
          dataQ_13 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_8095) begin
          dataQ_14 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_8131) begin
          dataQ_15 <= io_dataFromStorePorts_0;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_7574) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_7610) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_7646) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_7682) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_7718) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_7754) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_7790) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_7826) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_7862) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_7898) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_7934) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_7970) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_8006) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_8042) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_8078) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_8114) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_7591) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_7627) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_7663) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_7699) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_7735) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_7771) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_7807) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_7843) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_7879) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_7915) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_7951) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_7987) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_8023) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_8059) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_8095) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_8131) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1766;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1767;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1768;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1769;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1770;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1771;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1772;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1773;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1774;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1775;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1776;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1777;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1778;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1779;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1780;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1781;
    end
    if (reset) begin
      storeCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        storeCompleted_0 <= 1'h0;
      end else begin
        if (_T_3554) begin
          storeCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        storeCompleted_1 <= 1'h0;
      end else begin
        if (_T_3559) begin
          storeCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        storeCompleted_2 <= 1'h0;
      end else begin
        if (_T_3564) begin
          storeCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        storeCompleted_3 <= 1'h0;
      end else begin
        if (_T_3569) begin
          storeCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        storeCompleted_4 <= 1'h0;
      end else begin
        if (_T_3574) begin
          storeCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        storeCompleted_5 <= 1'h0;
      end else begin
        if (_T_3579) begin
          storeCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        storeCompleted_6 <= 1'h0;
      end else begin
        if (_T_3584) begin
          storeCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        storeCompleted_7 <= 1'h0;
      end else begin
        if (_T_3589) begin
          storeCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        storeCompleted_8 <= 1'h0;
      end else begin
        if (_T_3594) begin
          storeCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        storeCompleted_9 <= 1'h0;
      end else begin
        if (_T_3599) begin
          storeCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        storeCompleted_10 <= 1'h0;
      end else begin
        if (_T_3604) begin
          storeCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        storeCompleted_11 <= 1'h0;
      end else begin
        if (_T_3609) begin
          storeCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        storeCompleted_12 <= 1'h0;
      end else begin
        if (_T_3614) begin
          storeCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        storeCompleted_13 <= 1'h0;
      end else begin
        if (_T_3619) begin
          storeCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        storeCompleted_14 <= 1'h0;
      end else begin
        if (_T_3624) begin
          storeCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      storeCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        storeCompleted_15 <= 1'h0;
      end else begin
        if (_T_3629) begin
          storeCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2109;
      end else begin
        if (io_loadEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2113) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2121) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2139;
      end else begin
        if (io_loadEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2143) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2151) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2169;
      end else begin
        if (io_loadEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2173) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2181) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2199;
      end else begin
        if (io_loadEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2203) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2211) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2229;
      end else begin
        if (io_loadEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2233) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2241) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2259;
      end else begin
        if (io_loadEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2263) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2271) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2289;
      end else begin
        if (io_loadEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2293) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2301) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2319;
      end else begin
        if (io_loadEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2323) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2331) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2349;
      end else begin
        if (io_loadEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2353) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2361) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2379;
      end else begin
        if (io_loadEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2383) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2391) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2409;
      end else begin
        if (io_loadEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2413) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2421) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2439;
      end else begin
        if (io_loadEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2443) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2451) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2469;
      end else begin
        if (io_loadEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2473) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2481) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2499;
      end else begin
        if (io_loadEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2503) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2511) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2529;
      end else begin
        if (io_loadEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2533) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2541) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2559;
      end else begin
        if (io_loadEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2563) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2571) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousLoadHead <= io_loadHead;
  end
endmodule
module LOAD_QUEUE_LSQ_a( // @[:@4838.2]
  input         clock, // @[:@4839.4]
  input         reset, // @[:@4840.4]
  input         io_bbStart, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_0, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_1, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_2, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_3, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_4, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_5, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_6, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_7, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_8, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_9, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_10, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_11, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_12, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_13, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_14, // @[:@4841.4]
  input  [3:0]  io_bbLoadOffsets_15, // @[:@4841.4]
  input         io_bbNumLoads, // @[:@4841.4]
  output [3:0]  io_loadTail, // @[:@4841.4]
  output [3:0]  io_loadHead, // @[:@4841.4]
  output        io_loadEmpty, // @[:@4841.4]
  input  [3:0]  io_storeTail, // @[:@4841.4]
  input  [3:0]  io_storeHead, // @[:@4841.4]
  input         io_storeEmpty, // @[:@4841.4]
  input         io_storeAddrDone_0, // @[:@4841.4]
  input         io_storeAddrDone_1, // @[:@4841.4]
  input         io_storeAddrDone_2, // @[:@4841.4]
  input         io_storeAddrDone_3, // @[:@4841.4]
  input         io_storeAddrDone_4, // @[:@4841.4]
  input         io_storeAddrDone_5, // @[:@4841.4]
  input         io_storeAddrDone_6, // @[:@4841.4]
  input         io_storeAddrDone_7, // @[:@4841.4]
  input         io_storeAddrDone_8, // @[:@4841.4]
  input         io_storeAddrDone_9, // @[:@4841.4]
  input         io_storeAddrDone_10, // @[:@4841.4]
  input         io_storeAddrDone_11, // @[:@4841.4]
  input         io_storeAddrDone_12, // @[:@4841.4]
  input         io_storeAddrDone_13, // @[:@4841.4]
  input         io_storeAddrDone_14, // @[:@4841.4]
  input         io_storeAddrDone_15, // @[:@4841.4]
  input         io_storeDataDone_0, // @[:@4841.4]
  input         io_storeDataDone_1, // @[:@4841.4]
  input         io_storeDataDone_2, // @[:@4841.4]
  input         io_storeDataDone_3, // @[:@4841.4]
  input         io_storeDataDone_4, // @[:@4841.4]
  input         io_storeDataDone_5, // @[:@4841.4]
  input         io_storeDataDone_6, // @[:@4841.4]
  input         io_storeDataDone_7, // @[:@4841.4]
  input         io_storeDataDone_8, // @[:@4841.4]
  input         io_storeDataDone_9, // @[:@4841.4]
  input         io_storeDataDone_10, // @[:@4841.4]
  input         io_storeDataDone_11, // @[:@4841.4]
  input         io_storeDataDone_12, // @[:@4841.4]
  input         io_storeDataDone_13, // @[:@4841.4]
  input         io_storeDataDone_14, // @[:@4841.4]
  input         io_storeDataDone_15, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_0, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_1, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_2, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_3, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_4, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_5, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_6, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_7, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_8, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_9, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_10, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_11, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_12, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_13, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_14, // @[:@4841.4]
  input  [30:0] io_storeAddrQueue_15, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_0, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_1, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_2, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_3, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_4, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_5, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_6, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_7, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_8, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_9, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_10, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_11, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_12, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_13, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_14, // @[:@4841.4]
  input  [31:0] io_storeDataQueue_15, // @[:@4841.4]
  output        io_loadAddrDone_0, // @[:@4841.4]
  output        io_loadAddrDone_1, // @[:@4841.4]
  output        io_loadAddrDone_2, // @[:@4841.4]
  output        io_loadAddrDone_3, // @[:@4841.4]
  output        io_loadAddrDone_4, // @[:@4841.4]
  output        io_loadAddrDone_5, // @[:@4841.4]
  output        io_loadAddrDone_6, // @[:@4841.4]
  output        io_loadAddrDone_7, // @[:@4841.4]
  output        io_loadAddrDone_8, // @[:@4841.4]
  output        io_loadAddrDone_9, // @[:@4841.4]
  output        io_loadAddrDone_10, // @[:@4841.4]
  output        io_loadAddrDone_11, // @[:@4841.4]
  output        io_loadAddrDone_12, // @[:@4841.4]
  output        io_loadAddrDone_13, // @[:@4841.4]
  output        io_loadAddrDone_14, // @[:@4841.4]
  output        io_loadAddrDone_15, // @[:@4841.4]
  output        io_loadDataDone_0, // @[:@4841.4]
  output        io_loadDataDone_1, // @[:@4841.4]
  output        io_loadDataDone_2, // @[:@4841.4]
  output        io_loadDataDone_3, // @[:@4841.4]
  output        io_loadDataDone_4, // @[:@4841.4]
  output        io_loadDataDone_5, // @[:@4841.4]
  output        io_loadDataDone_6, // @[:@4841.4]
  output        io_loadDataDone_7, // @[:@4841.4]
  output        io_loadDataDone_8, // @[:@4841.4]
  output        io_loadDataDone_9, // @[:@4841.4]
  output        io_loadDataDone_10, // @[:@4841.4]
  output        io_loadDataDone_11, // @[:@4841.4]
  output        io_loadDataDone_12, // @[:@4841.4]
  output        io_loadDataDone_13, // @[:@4841.4]
  output        io_loadDataDone_14, // @[:@4841.4]
  output        io_loadDataDone_15, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_0, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_1, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_2, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_3, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_4, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_5, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_6, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_7, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_8, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_9, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_10, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_11, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_12, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_13, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_14, // @[:@4841.4]
  output [30:0] io_loadAddrQueue_15, // @[:@4841.4]
  input         io_loadAddrEnable_0, // @[:@4841.4]
  input  [30:0] io_addrFromLoadPorts_0, // @[:@4841.4]
  input         io_loadPorts_0_ready, // @[:@4841.4]
  output        io_loadPorts_0_valid, // @[:@4841.4]
  output [31:0] io_loadPorts_0_bits, // @[:@4841.4]
  input  [31:0] io_loadDataFromMem, // @[:@4841.4]
  output [30:0] io_loadAddrToMem, // @[:@4841.4]
  input  [31:0] io_loadQIdxForDataIn, // @[:@4841.4]
  input         io_loadQIdxForDataInValid, // @[:@4841.4]
  input         io_loadQIdxForAddrOut_ready, // @[:@4841.4]
  output        io_loadQIdxForAddrOut_valid, // @[:@4841.4]
  output [3:0]  io_loadQIdxForAddrOut_bits // @[:@4841.4]
);
  reg [3:0] head; // @[AxiLoadQueue.scala 50:21:@4843.4]
  reg [31:0] _RAND_0;
  reg [3:0] tail; // @[AxiLoadQueue.scala 51:21:@4844.4]
  reg [31:0] _RAND_1;
  reg [3:0] offsetQ_0; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_2;
  reg [3:0] offsetQ_1; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_3;
  reg [3:0] offsetQ_2; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_4;
  reg [3:0] offsetQ_3; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_5;
  reg [3:0] offsetQ_4; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_6;
  reg [3:0] offsetQ_5; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_7;
  reg [3:0] offsetQ_6; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_8;
  reg [3:0] offsetQ_7; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_9;
  reg [3:0] offsetQ_8; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_10;
  reg [3:0] offsetQ_9; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_11;
  reg [3:0] offsetQ_10; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_12;
  reg [3:0] offsetQ_11; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_13;
  reg [3:0] offsetQ_12; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_14;
  reg [3:0] offsetQ_13; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_15;
  reg [3:0] offsetQ_14; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_16;
  reg [3:0] offsetQ_15; // @[AxiLoadQueue.scala 53:24:@4862.4]
  reg [31:0] _RAND_17;
  reg  portQ_0; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_18;
  reg  portQ_1; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_19;
  reg  portQ_2; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_20;
  reg  portQ_3; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_21;
  reg  portQ_4; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_22;
  reg  portQ_5; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_23;
  reg  portQ_6; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_24;
  reg  portQ_7; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_25;
  reg  portQ_8; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_26;
  reg  portQ_9; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_27;
  reg  portQ_10; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_28;
  reg  portQ_11; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_29;
  reg  portQ_12; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_30;
  reg  portQ_13; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_31;
  reg  portQ_14; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_32;
  reg  portQ_15; // @[AxiLoadQueue.scala 54:22:@4880.4]
  reg [31:0] _RAND_33;
  reg [30:0] addrQ_0; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_34;
  reg [30:0] addrQ_1; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_35;
  reg [30:0] addrQ_2; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_36;
  reg [30:0] addrQ_3; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_37;
  reg [30:0] addrQ_4; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_38;
  reg [30:0] addrQ_5; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_39;
  reg [30:0] addrQ_6; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_40;
  reg [30:0] addrQ_7; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_41;
  reg [30:0] addrQ_8; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_42;
  reg [30:0] addrQ_9; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_43;
  reg [30:0] addrQ_10; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_44;
  reg [30:0] addrQ_11; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_45;
  reg [30:0] addrQ_12; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_46;
  reg [30:0] addrQ_13; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_47;
  reg [30:0] addrQ_14; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_48;
  reg [30:0] addrQ_15; // @[AxiLoadQueue.scala 55:22:@4898.4]
  reg [31:0] _RAND_49;
  reg [31:0] dataQ_0; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_50;
  reg [31:0] dataQ_1; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_51;
  reg [31:0] dataQ_2; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_52;
  reg [31:0] dataQ_3; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_53;
  reg [31:0] dataQ_4; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_54;
  reg [31:0] dataQ_5; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_55;
  reg [31:0] dataQ_6; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_56;
  reg [31:0] dataQ_7; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_57;
  reg [31:0] dataQ_8; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_58;
  reg [31:0] dataQ_9; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_59;
  reg [31:0] dataQ_10; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_60;
  reg [31:0] dataQ_11; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_61;
  reg [31:0] dataQ_12; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_62;
  reg [31:0] dataQ_13; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_63;
  reg [31:0] dataQ_14; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_64;
  reg [31:0] dataQ_15; // @[AxiLoadQueue.scala 56:22:@4916.4]
  reg [31:0] _RAND_65;
  reg  addrKnown_0; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_66;
  reg  addrKnown_1; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_67;
  reg  addrKnown_2; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_68;
  reg  addrKnown_3; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_69;
  reg  addrKnown_4; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_70;
  reg  addrKnown_5; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_71;
  reg  addrKnown_6; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_72;
  reg  addrKnown_7; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_73;
  reg  addrKnown_8; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_74;
  reg  addrKnown_9; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_75;
  reg  addrKnown_10; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_76;
  reg  addrKnown_11; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_77;
  reg  addrKnown_12; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_78;
  reg  addrKnown_13; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_79;
  reg  addrKnown_14; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_80;
  reg  addrKnown_15; // @[AxiLoadQueue.scala 57:26:@4934.4]
  reg [31:0] _RAND_81;
  reg  dataKnown_0; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_82;
  reg  dataKnown_1; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_83;
  reg  dataKnown_2; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_84;
  reg  dataKnown_3; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_85;
  reg  dataKnown_4; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_86;
  reg  dataKnown_5; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_87;
  reg  dataKnown_6; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_88;
  reg  dataKnown_7; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_89;
  reg  dataKnown_8; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_90;
  reg  dataKnown_9; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_91;
  reg  dataKnown_10; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_92;
  reg  dataKnown_11; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_93;
  reg  dataKnown_12; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_94;
  reg  dataKnown_13; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_95;
  reg  dataKnown_14; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_96;
  reg  dataKnown_15; // @[AxiLoadQueue.scala 58:26:@4952.4]
  reg [31:0] _RAND_97;
  reg  loadCompleted_0; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_98;
  reg  loadCompleted_1; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_99;
  reg  loadCompleted_2; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_100;
  reg  loadCompleted_3; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_101;
  reg  loadCompleted_4; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_102;
  reg  loadCompleted_5; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_103;
  reg  loadCompleted_6; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_104;
  reg  loadCompleted_7; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_105;
  reg  loadCompleted_8; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_106;
  reg  loadCompleted_9; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_107;
  reg  loadCompleted_10; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_108;
  reg  loadCompleted_11; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_109;
  reg  loadCompleted_12; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_110;
  reg  loadCompleted_13; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_111;
  reg  loadCompleted_14; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_112;
  reg  loadCompleted_15; // @[AxiLoadQueue.scala 59:30:@4970.4]
  reg [31:0] _RAND_113;
  reg  allocatedEntries_0; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_114;
  reg  allocatedEntries_1; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_115;
  reg  allocatedEntries_2; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_116;
  reg  allocatedEntries_3; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_117;
  reg  allocatedEntries_4; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_118;
  reg  allocatedEntries_5; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_119;
  reg  allocatedEntries_6; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_120;
  reg  allocatedEntries_7; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_121;
  reg  allocatedEntries_8; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_122;
  reg  allocatedEntries_9; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_123;
  reg  allocatedEntries_10; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_124;
  reg  allocatedEntries_11; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_125;
  reg  allocatedEntries_12; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_126;
  reg  allocatedEntries_13; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_127;
  reg  allocatedEntries_14; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_128;
  reg  allocatedEntries_15; // @[AxiLoadQueue.scala 60:33:@4988.4]
  reg [31:0] _RAND_129;
  reg  bypassInitiated_0; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_130;
  reg  bypassInitiated_1; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_131;
  reg  bypassInitiated_2; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_132;
  reg  bypassInitiated_3; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_133;
  reg  bypassInitiated_4; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_134;
  reg  bypassInitiated_5; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_135;
  reg  bypassInitiated_6; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_136;
  reg  bypassInitiated_7; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_137;
  reg  bypassInitiated_8; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_138;
  reg  bypassInitiated_9; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_139;
  reg  bypassInitiated_10; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_140;
  reg  bypassInitiated_11; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_141;
  reg  bypassInitiated_12; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_142;
  reg  bypassInitiated_13; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_143;
  reg  bypassInitiated_14; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_144;
  reg  bypassInitiated_15; // @[AxiLoadQueue.scala 61:32:@5006.4]
  reg [31:0] _RAND_145;
  reg  checkBits_0; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_146;
  reg  checkBits_1; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_147;
  reg  checkBits_2; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_148;
  reg  checkBits_3; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_149;
  reg  checkBits_4; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_150;
  reg  checkBits_5; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_151;
  reg  checkBits_6; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_152;
  reg  checkBits_7; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_153;
  reg  checkBits_8; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_154;
  reg  checkBits_9; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_155;
  reg  checkBits_10; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_156;
  reg  checkBits_11; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_157;
  reg  checkBits_12; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_158;
  reg  checkBits_13; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_159;
  reg  checkBits_14; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_160;
  reg  checkBits_15; // @[AxiLoadQueue.scala 62:26:@5024.4]
  reg [31:0] _RAND_161;
  wire [5:0] _GEN_2276; // @[util.scala 14:20:@5026.4]
  wire [6:0] _T_1722; // @[util.scala 14:20:@5026.4]
  wire [6:0] _T_1723; // @[util.scala 14:20:@5027.4]
  wire [5:0] _T_1724; // @[util.scala 14:20:@5028.4]
  wire [5:0] _GEN_0; // @[util.scala 14:25:@5029.4]
  wire [4:0] _T_1725; // @[util.scala 14:25:@5029.4]
  wire [4:0] _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5030.4]
  wire  _T_1726; // @[AxiLoadQueue.scala 71:46:@5030.4]
  wire  initBits_0; // @[AxiLoadQueue.scala 71:63:@5031.4]
  wire [6:0] _T_1731; // @[util.scala 14:20:@5033.4]
  wire [6:0] _T_1732; // @[util.scala 14:20:@5034.4]
  wire [5:0] _T_1733; // @[util.scala 14:20:@5035.4]
  wire [5:0] _GEN_16; // @[util.scala 14:25:@5036.4]
  wire [4:0] _T_1734; // @[util.scala 14:25:@5036.4]
  wire  _T_1735; // @[AxiLoadQueue.scala 71:46:@5037.4]
  wire  initBits_1; // @[AxiLoadQueue.scala 71:63:@5038.4]
  wire [6:0] _T_1740; // @[util.scala 14:20:@5040.4]
  wire [6:0] _T_1741; // @[util.scala 14:20:@5041.4]
  wire [5:0] _T_1742; // @[util.scala 14:20:@5042.4]
  wire [5:0] _GEN_17; // @[util.scala 14:25:@5043.4]
  wire [4:0] _T_1743; // @[util.scala 14:25:@5043.4]
  wire  _T_1744; // @[AxiLoadQueue.scala 71:46:@5044.4]
  wire  initBits_2; // @[AxiLoadQueue.scala 71:63:@5045.4]
  wire [6:0] _T_1749; // @[util.scala 14:20:@5047.4]
  wire [6:0] _T_1750; // @[util.scala 14:20:@5048.4]
  wire [5:0] _T_1751; // @[util.scala 14:20:@5049.4]
  wire [5:0] _GEN_18; // @[util.scala 14:25:@5050.4]
  wire [4:0] _T_1752; // @[util.scala 14:25:@5050.4]
  wire  _T_1753; // @[AxiLoadQueue.scala 71:46:@5051.4]
  wire  initBits_3; // @[AxiLoadQueue.scala 71:63:@5052.4]
  wire [6:0] _T_1758; // @[util.scala 14:20:@5054.4]
  wire [6:0] _T_1759; // @[util.scala 14:20:@5055.4]
  wire [5:0] _T_1760; // @[util.scala 14:20:@5056.4]
  wire [5:0] _GEN_19; // @[util.scala 14:25:@5057.4]
  wire [4:0] _T_1761; // @[util.scala 14:25:@5057.4]
  wire  _T_1762; // @[AxiLoadQueue.scala 71:46:@5058.4]
  wire  initBits_4; // @[AxiLoadQueue.scala 71:63:@5059.4]
  wire [6:0] _T_1767; // @[util.scala 14:20:@5061.4]
  wire [6:0] _T_1768; // @[util.scala 14:20:@5062.4]
  wire [5:0] _T_1769; // @[util.scala 14:20:@5063.4]
  wire [5:0] _GEN_20; // @[util.scala 14:25:@5064.4]
  wire [4:0] _T_1770; // @[util.scala 14:25:@5064.4]
  wire  _T_1771; // @[AxiLoadQueue.scala 71:46:@5065.4]
  wire  initBits_5; // @[AxiLoadQueue.scala 71:63:@5066.4]
  wire [6:0] _T_1776; // @[util.scala 14:20:@5068.4]
  wire [6:0] _T_1777; // @[util.scala 14:20:@5069.4]
  wire [5:0] _T_1778; // @[util.scala 14:20:@5070.4]
  wire [5:0] _GEN_21; // @[util.scala 14:25:@5071.4]
  wire [4:0] _T_1779; // @[util.scala 14:25:@5071.4]
  wire  _T_1780; // @[AxiLoadQueue.scala 71:46:@5072.4]
  wire  initBits_6; // @[AxiLoadQueue.scala 71:63:@5073.4]
  wire [6:0] _T_1785; // @[util.scala 14:20:@5075.4]
  wire [6:0] _T_1786; // @[util.scala 14:20:@5076.4]
  wire [5:0] _T_1787; // @[util.scala 14:20:@5077.4]
  wire [5:0] _GEN_22; // @[util.scala 14:25:@5078.4]
  wire [4:0] _T_1788; // @[util.scala 14:25:@5078.4]
  wire  _T_1789; // @[AxiLoadQueue.scala 71:46:@5079.4]
  wire  initBits_7; // @[AxiLoadQueue.scala 71:63:@5080.4]
  wire [6:0] _T_1794; // @[util.scala 14:20:@5082.4]
  wire [6:0] _T_1795; // @[util.scala 14:20:@5083.4]
  wire [5:0] _T_1796; // @[util.scala 14:20:@5084.4]
  wire [5:0] _GEN_23; // @[util.scala 14:25:@5085.4]
  wire [4:0] _T_1797; // @[util.scala 14:25:@5085.4]
  wire  _T_1798; // @[AxiLoadQueue.scala 71:46:@5086.4]
  wire  initBits_8; // @[AxiLoadQueue.scala 71:63:@5087.4]
  wire [6:0] _T_1803; // @[util.scala 14:20:@5089.4]
  wire [6:0] _T_1804; // @[util.scala 14:20:@5090.4]
  wire [5:0] _T_1805; // @[util.scala 14:20:@5091.4]
  wire [5:0] _GEN_24; // @[util.scala 14:25:@5092.4]
  wire [4:0] _T_1806; // @[util.scala 14:25:@5092.4]
  wire  _T_1807; // @[AxiLoadQueue.scala 71:46:@5093.4]
  wire  initBits_9; // @[AxiLoadQueue.scala 71:63:@5094.4]
  wire [6:0] _T_1812; // @[util.scala 14:20:@5096.4]
  wire [6:0] _T_1813; // @[util.scala 14:20:@5097.4]
  wire [5:0] _T_1814; // @[util.scala 14:20:@5098.4]
  wire [5:0] _GEN_25; // @[util.scala 14:25:@5099.4]
  wire [4:0] _T_1815; // @[util.scala 14:25:@5099.4]
  wire  _T_1816; // @[AxiLoadQueue.scala 71:46:@5100.4]
  wire  initBits_10; // @[AxiLoadQueue.scala 71:63:@5101.4]
  wire [6:0] _T_1821; // @[util.scala 14:20:@5103.4]
  wire [6:0] _T_1822; // @[util.scala 14:20:@5104.4]
  wire [5:0] _T_1823; // @[util.scala 14:20:@5105.4]
  wire [5:0] _GEN_26; // @[util.scala 14:25:@5106.4]
  wire [4:0] _T_1824; // @[util.scala 14:25:@5106.4]
  wire  _T_1825; // @[AxiLoadQueue.scala 71:46:@5107.4]
  wire  initBits_11; // @[AxiLoadQueue.scala 71:63:@5108.4]
  wire [6:0] _T_1830; // @[util.scala 14:20:@5110.4]
  wire [6:0] _T_1831; // @[util.scala 14:20:@5111.4]
  wire [5:0] _T_1832; // @[util.scala 14:20:@5112.4]
  wire [5:0] _GEN_27; // @[util.scala 14:25:@5113.4]
  wire [4:0] _T_1833; // @[util.scala 14:25:@5113.4]
  wire  _T_1834; // @[AxiLoadQueue.scala 71:46:@5114.4]
  wire  initBits_12; // @[AxiLoadQueue.scala 71:63:@5115.4]
  wire [6:0] _T_1839; // @[util.scala 14:20:@5117.4]
  wire [6:0] _T_1840; // @[util.scala 14:20:@5118.4]
  wire [5:0] _T_1841; // @[util.scala 14:20:@5119.4]
  wire [5:0] _GEN_28; // @[util.scala 14:25:@5120.4]
  wire [4:0] _T_1842; // @[util.scala 14:25:@5120.4]
  wire  _T_1843; // @[AxiLoadQueue.scala 71:46:@5121.4]
  wire  initBits_13; // @[AxiLoadQueue.scala 71:63:@5122.4]
  wire [6:0] _T_1848; // @[util.scala 14:20:@5124.4]
  wire [6:0] _T_1849; // @[util.scala 14:20:@5125.4]
  wire [5:0] _T_1850; // @[util.scala 14:20:@5126.4]
  wire [5:0] _GEN_29; // @[util.scala 14:25:@5127.4]
  wire [4:0] _T_1851; // @[util.scala 14:25:@5127.4]
  wire  _T_1852; // @[AxiLoadQueue.scala 71:46:@5128.4]
  wire  initBits_14; // @[AxiLoadQueue.scala 71:63:@5129.4]
  wire [6:0] _T_1857; // @[util.scala 14:20:@5131.4]
  wire [6:0] _T_1858; // @[util.scala 14:20:@5132.4]
  wire [5:0] _T_1859; // @[util.scala 14:20:@5133.4]
  wire [5:0] _GEN_30; // @[util.scala 14:25:@5134.4]
  wire [4:0] _T_1860; // @[util.scala 14:25:@5134.4]
  wire  _T_1861; // @[AxiLoadQueue.scala 71:46:@5135.4]
  wire  initBits_15; // @[AxiLoadQueue.scala 71:63:@5136.4]
  wire  _T_1884; // @[AxiLoadQueue.scala 73:78:@5154.4]
  wire  _T_1885; // @[AxiLoadQueue.scala 73:78:@5155.4]
  wire  _T_1886; // @[AxiLoadQueue.scala 73:78:@5156.4]
  wire  _T_1887; // @[AxiLoadQueue.scala 73:78:@5157.4]
  wire  _T_1888; // @[AxiLoadQueue.scala 73:78:@5158.4]
  wire  _T_1889; // @[AxiLoadQueue.scala 73:78:@5159.4]
  wire  _T_1890; // @[AxiLoadQueue.scala 73:78:@5160.4]
  wire  _T_1891; // @[AxiLoadQueue.scala 73:78:@5161.4]
  wire  _T_1892; // @[AxiLoadQueue.scala 73:78:@5162.4]
  wire  _T_1893; // @[AxiLoadQueue.scala 73:78:@5163.4]
  wire  _T_1894; // @[AxiLoadQueue.scala 73:78:@5164.4]
  wire  _T_1895; // @[AxiLoadQueue.scala 73:78:@5165.4]
  wire  _T_1896; // @[AxiLoadQueue.scala 73:78:@5166.4]
  wire  _T_1897; // @[AxiLoadQueue.scala 73:78:@5167.4]
  wire  _T_1898; // @[AxiLoadQueue.scala 73:78:@5168.4]
  wire  _T_1899; // @[AxiLoadQueue.scala 73:78:@5169.4]
  wire [3:0] _T_1930; // @[:@5209.6]
  wire [3:0] _GEN_1; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_2; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_3; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_4; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_5; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_6; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_7; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_8; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_9; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_10; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_11; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_12; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_13; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_14; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_15; // @[AxiLoadQueue.scala 77:20:@5210.6]
  wire [3:0] _GEN_32; // @[AxiLoadQueue.scala 76:25:@5203.4]
  wire  _GEN_33; // @[AxiLoadQueue.scala 76:25:@5203.4]
  wire [3:0] _T_1948; // @[:@5225.6]
  wire [3:0] _GEN_35; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_36; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_37; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_38; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_39; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_40; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_41; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_42; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_43; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_44; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_45; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_46; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_47; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_48; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_49; // @[AxiLoadQueue.scala 77:20:@5226.6]
  wire [3:0] _GEN_66; // @[AxiLoadQueue.scala 76:25:@5219.4]
  wire  _GEN_67; // @[AxiLoadQueue.scala 76:25:@5219.4]
  wire [3:0] _T_1966; // @[:@5241.6]
  wire [3:0] _GEN_69; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_70; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_71; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_72; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_73; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_74; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_75; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_76; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_77; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_78; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_79; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_80; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_81; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_82; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_83; // @[AxiLoadQueue.scala 77:20:@5242.6]
  wire [3:0] _GEN_100; // @[AxiLoadQueue.scala 76:25:@5235.4]
  wire  _GEN_101; // @[AxiLoadQueue.scala 76:25:@5235.4]
  wire [3:0] _T_1984; // @[:@5257.6]
  wire [3:0] _GEN_103; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_104; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_105; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_106; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_107; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_108; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_109; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_110; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_111; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_112; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_113; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_114; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_115; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_116; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_117; // @[AxiLoadQueue.scala 77:20:@5258.6]
  wire [3:0] _GEN_134; // @[AxiLoadQueue.scala 76:25:@5251.4]
  wire  _GEN_135; // @[AxiLoadQueue.scala 76:25:@5251.4]
  wire [3:0] _T_2002; // @[:@5273.6]
  wire [3:0] _GEN_137; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_138; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_139; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_140; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_141; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_142; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_143; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_144; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_145; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_146; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_147; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_148; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_149; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_150; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_151; // @[AxiLoadQueue.scala 77:20:@5274.6]
  wire [3:0] _GEN_168; // @[AxiLoadQueue.scala 76:25:@5267.4]
  wire  _GEN_169; // @[AxiLoadQueue.scala 76:25:@5267.4]
  wire [3:0] _T_2020; // @[:@5289.6]
  wire [3:0] _GEN_171; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_172; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_173; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_174; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_175; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_176; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_177; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_178; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_179; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_180; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_181; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_182; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_183; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_184; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_185; // @[AxiLoadQueue.scala 77:20:@5290.6]
  wire [3:0] _GEN_202; // @[AxiLoadQueue.scala 76:25:@5283.4]
  wire  _GEN_203; // @[AxiLoadQueue.scala 76:25:@5283.4]
  wire [3:0] _T_2038; // @[:@5305.6]
  wire [3:0] _GEN_205; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_206; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_207; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_208; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_209; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_210; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_211; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_212; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_213; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_214; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_215; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_216; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_217; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_218; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_219; // @[AxiLoadQueue.scala 77:20:@5306.6]
  wire [3:0] _GEN_236; // @[AxiLoadQueue.scala 76:25:@5299.4]
  wire  _GEN_237; // @[AxiLoadQueue.scala 76:25:@5299.4]
  wire [3:0] _T_2056; // @[:@5321.6]
  wire [3:0] _GEN_239; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_240; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_241; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_242; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_243; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_244; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_245; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_246; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_247; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_248; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_249; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_250; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_251; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_252; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_253; // @[AxiLoadQueue.scala 77:20:@5322.6]
  wire [3:0] _GEN_270; // @[AxiLoadQueue.scala 76:25:@5315.4]
  wire  _GEN_271; // @[AxiLoadQueue.scala 76:25:@5315.4]
  wire [3:0] _T_2074; // @[:@5337.6]
  wire [3:0] _GEN_273; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_274; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_275; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_276; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_277; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_278; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_279; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_280; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_281; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_282; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_283; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_284; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_285; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_286; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_287; // @[AxiLoadQueue.scala 77:20:@5338.6]
  wire [3:0] _GEN_304; // @[AxiLoadQueue.scala 76:25:@5331.4]
  wire  _GEN_305; // @[AxiLoadQueue.scala 76:25:@5331.4]
  wire [3:0] _T_2092; // @[:@5353.6]
  wire [3:0] _GEN_307; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_308; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_309; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_310; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_311; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_312; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_313; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_314; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_315; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_316; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_317; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_318; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_319; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_320; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_321; // @[AxiLoadQueue.scala 77:20:@5354.6]
  wire [3:0] _GEN_338; // @[AxiLoadQueue.scala 76:25:@5347.4]
  wire  _GEN_339; // @[AxiLoadQueue.scala 76:25:@5347.4]
  wire [3:0] _T_2110; // @[:@5369.6]
  wire [3:0] _GEN_341; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_342; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_343; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_344; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_345; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_346; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_347; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_348; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_349; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_350; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_351; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_352; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_353; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_354; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_355; // @[AxiLoadQueue.scala 77:20:@5370.6]
  wire [3:0] _GEN_372; // @[AxiLoadQueue.scala 76:25:@5363.4]
  wire  _GEN_373; // @[AxiLoadQueue.scala 76:25:@5363.4]
  wire [3:0] _T_2128; // @[:@5385.6]
  wire [3:0] _GEN_375; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_376; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_377; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_378; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_379; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_380; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_381; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_382; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_383; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_384; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_385; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_386; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_387; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_388; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_389; // @[AxiLoadQueue.scala 77:20:@5386.6]
  wire [3:0] _GEN_406; // @[AxiLoadQueue.scala 76:25:@5379.4]
  wire  _GEN_407; // @[AxiLoadQueue.scala 76:25:@5379.4]
  wire [3:0] _T_2146; // @[:@5401.6]
  wire [3:0] _GEN_409; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_410; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_411; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_412; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_413; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_414; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_415; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_416; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_417; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_418; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_419; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_420; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_421; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_422; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_423; // @[AxiLoadQueue.scala 77:20:@5402.6]
  wire [3:0] _GEN_440; // @[AxiLoadQueue.scala 76:25:@5395.4]
  wire  _GEN_441; // @[AxiLoadQueue.scala 76:25:@5395.4]
  wire [3:0] _T_2164; // @[:@5417.6]
  wire [3:0] _GEN_443; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_444; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_445; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_446; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_447; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_448; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_449; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_450; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_451; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_452; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_453; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_454; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_455; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_456; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_457; // @[AxiLoadQueue.scala 77:20:@5418.6]
  wire [3:0] _GEN_474; // @[AxiLoadQueue.scala 76:25:@5411.4]
  wire  _GEN_475; // @[AxiLoadQueue.scala 76:25:@5411.4]
  wire [3:0] _T_2182; // @[:@5433.6]
  wire [3:0] _GEN_477; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_478; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_479; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_480; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_481; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_482; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_483; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_484; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_485; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_486; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_487; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_488; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_489; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_490; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_491; // @[AxiLoadQueue.scala 77:20:@5434.6]
  wire [3:0] _GEN_508; // @[AxiLoadQueue.scala 76:25:@5427.4]
  wire  _GEN_509; // @[AxiLoadQueue.scala 76:25:@5427.4]
  wire [3:0] _T_2200; // @[:@5449.6]
  wire [3:0] _GEN_511; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_512; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_513; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_514; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_515; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_516; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_517; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_518; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_519; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_520; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_521; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_522; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_523; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_524; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_525; // @[AxiLoadQueue.scala 77:20:@5450.6]
  wire [3:0] _GEN_542; // @[AxiLoadQueue.scala 76:25:@5443.4]
  wire  _GEN_543; // @[AxiLoadQueue.scala 76:25:@5443.4]
  reg [3:0] previousStoreHead; // @[AxiLoadQueue.scala 93:34:@5459.4]
  reg [31:0] _RAND_162;
  wire [4:0] _T_2222; // @[util.scala 10:8:@5468.6]
  wire [4:0] _GEN_31; // @[util.scala 10:14:@5469.6]
  wire [4:0] _T_2223; // @[util.scala 10:14:@5469.6]
  wire [4:0] _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5470.6]
  wire  _T_2224; // @[AxiLoadQueue.scala 97:56:@5470.6]
  wire  _T_2225; // @[AxiLoadQueue.scala 96:50:@5471.6]
  wire  _T_2227; // @[AxiLoadQueue.scala 96:34:@5472.6]
  wire  _T_2229; // @[AxiLoadQueue.scala 101:36:@5480.8]
  wire  _T_2230; // @[AxiLoadQueue.scala 101:86:@5481.8]
  wire  _T_2231; // @[AxiLoadQueue.scala 101:61:@5482.8]
  wire  _T_2233; // @[AxiLoadQueue.scala 103:36:@5487.10]
  wire  _T_2234; // @[AxiLoadQueue.scala 103:69:@5488.10]
  wire  _T_2235; // @[AxiLoadQueue.scala 104:31:@5489.10]
  wire  _T_2236; // @[AxiLoadQueue.scala 103:94:@5490.10]
  wire  _T_2238; // @[AxiLoadQueue.scala 103:54:@5491.10]
  wire  _T_2239; // @[AxiLoadQueue.scala 103:51:@5492.10]
  wire  _GEN_560; // @[AxiLoadQueue.scala 104:53:@5493.10]
  wire  _GEN_561; // @[AxiLoadQueue.scala 101:102:@5483.8]
  wire  _GEN_562; // @[AxiLoadQueue.scala 99:27:@5476.6]
  wire  _GEN_563; // @[AxiLoadQueue.scala 95:34:@5461.4]
  wire [4:0] _T_2252; // @[util.scala 10:8:@5504.6]
  wire [4:0] _GEN_34; // @[util.scala 10:14:@5505.6]
  wire [4:0] _T_2253; // @[util.scala 10:14:@5505.6]
  wire  _T_2254; // @[AxiLoadQueue.scala 97:56:@5506.6]
  wire  _T_2255; // @[AxiLoadQueue.scala 96:50:@5507.6]
  wire  _T_2257; // @[AxiLoadQueue.scala 96:34:@5508.6]
  wire  _T_2259; // @[AxiLoadQueue.scala 101:36:@5516.8]
  wire  _T_2260; // @[AxiLoadQueue.scala 101:86:@5517.8]
  wire  _T_2261; // @[AxiLoadQueue.scala 101:61:@5518.8]
  wire  _T_2264; // @[AxiLoadQueue.scala 103:69:@5524.10]
  wire  _T_2265; // @[AxiLoadQueue.scala 104:31:@5525.10]
  wire  _T_2266; // @[AxiLoadQueue.scala 103:94:@5526.10]
  wire  _T_2268; // @[AxiLoadQueue.scala 103:54:@5527.10]
  wire  _T_2269; // @[AxiLoadQueue.scala 103:51:@5528.10]
  wire  _GEN_580; // @[AxiLoadQueue.scala 104:53:@5529.10]
  wire  _GEN_581; // @[AxiLoadQueue.scala 101:102:@5519.8]
  wire  _GEN_582; // @[AxiLoadQueue.scala 99:27:@5512.6]
  wire  _GEN_583; // @[AxiLoadQueue.scala 95:34:@5497.4]
  wire [4:0] _T_2282; // @[util.scala 10:8:@5540.6]
  wire [4:0] _GEN_50; // @[util.scala 10:14:@5541.6]
  wire [4:0] _T_2283; // @[util.scala 10:14:@5541.6]
  wire  _T_2284; // @[AxiLoadQueue.scala 97:56:@5542.6]
  wire  _T_2285; // @[AxiLoadQueue.scala 96:50:@5543.6]
  wire  _T_2287; // @[AxiLoadQueue.scala 96:34:@5544.6]
  wire  _T_2289; // @[AxiLoadQueue.scala 101:36:@5552.8]
  wire  _T_2290; // @[AxiLoadQueue.scala 101:86:@5553.8]
  wire  _T_2291; // @[AxiLoadQueue.scala 101:61:@5554.8]
  wire  _T_2294; // @[AxiLoadQueue.scala 103:69:@5560.10]
  wire  _T_2295; // @[AxiLoadQueue.scala 104:31:@5561.10]
  wire  _T_2296; // @[AxiLoadQueue.scala 103:94:@5562.10]
  wire  _T_2298; // @[AxiLoadQueue.scala 103:54:@5563.10]
  wire  _T_2299; // @[AxiLoadQueue.scala 103:51:@5564.10]
  wire  _GEN_600; // @[AxiLoadQueue.scala 104:53:@5565.10]
  wire  _GEN_601; // @[AxiLoadQueue.scala 101:102:@5555.8]
  wire  _GEN_602; // @[AxiLoadQueue.scala 99:27:@5548.6]
  wire  _GEN_603; // @[AxiLoadQueue.scala 95:34:@5533.4]
  wire [4:0] _T_2312; // @[util.scala 10:8:@5576.6]
  wire [4:0] _GEN_51; // @[util.scala 10:14:@5577.6]
  wire [4:0] _T_2313; // @[util.scala 10:14:@5577.6]
  wire  _T_2314; // @[AxiLoadQueue.scala 97:56:@5578.6]
  wire  _T_2315; // @[AxiLoadQueue.scala 96:50:@5579.6]
  wire  _T_2317; // @[AxiLoadQueue.scala 96:34:@5580.6]
  wire  _T_2319; // @[AxiLoadQueue.scala 101:36:@5588.8]
  wire  _T_2320; // @[AxiLoadQueue.scala 101:86:@5589.8]
  wire  _T_2321; // @[AxiLoadQueue.scala 101:61:@5590.8]
  wire  _T_2324; // @[AxiLoadQueue.scala 103:69:@5596.10]
  wire  _T_2325; // @[AxiLoadQueue.scala 104:31:@5597.10]
  wire  _T_2326; // @[AxiLoadQueue.scala 103:94:@5598.10]
  wire  _T_2328; // @[AxiLoadQueue.scala 103:54:@5599.10]
  wire  _T_2329; // @[AxiLoadQueue.scala 103:51:@5600.10]
  wire  _GEN_620; // @[AxiLoadQueue.scala 104:53:@5601.10]
  wire  _GEN_621; // @[AxiLoadQueue.scala 101:102:@5591.8]
  wire  _GEN_622; // @[AxiLoadQueue.scala 99:27:@5584.6]
  wire  _GEN_623; // @[AxiLoadQueue.scala 95:34:@5569.4]
  wire [4:0] _T_2342; // @[util.scala 10:8:@5612.6]
  wire [4:0] _GEN_52; // @[util.scala 10:14:@5613.6]
  wire [4:0] _T_2343; // @[util.scala 10:14:@5613.6]
  wire  _T_2344; // @[AxiLoadQueue.scala 97:56:@5614.6]
  wire  _T_2345; // @[AxiLoadQueue.scala 96:50:@5615.6]
  wire  _T_2347; // @[AxiLoadQueue.scala 96:34:@5616.6]
  wire  _T_2349; // @[AxiLoadQueue.scala 101:36:@5624.8]
  wire  _T_2350; // @[AxiLoadQueue.scala 101:86:@5625.8]
  wire  _T_2351; // @[AxiLoadQueue.scala 101:61:@5626.8]
  wire  _T_2354; // @[AxiLoadQueue.scala 103:69:@5632.10]
  wire  _T_2355; // @[AxiLoadQueue.scala 104:31:@5633.10]
  wire  _T_2356; // @[AxiLoadQueue.scala 103:94:@5634.10]
  wire  _T_2358; // @[AxiLoadQueue.scala 103:54:@5635.10]
  wire  _T_2359; // @[AxiLoadQueue.scala 103:51:@5636.10]
  wire  _GEN_640; // @[AxiLoadQueue.scala 104:53:@5637.10]
  wire  _GEN_641; // @[AxiLoadQueue.scala 101:102:@5627.8]
  wire  _GEN_642; // @[AxiLoadQueue.scala 99:27:@5620.6]
  wire  _GEN_643; // @[AxiLoadQueue.scala 95:34:@5605.4]
  wire [4:0] _T_2372; // @[util.scala 10:8:@5648.6]
  wire [4:0] _GEN_53; // @[util.scala 10:14:@5649.6]
  wire [4:0] _T_2373; // @[util.scala 10:14:@5649.6]
  wire  _T_2374; // @[AxiLoadQueue.scala 97:56:@5650.6]
  wire  _T_2375; // @[AxiLoadQueue.scala 96:50:@5651.6]
  wire  _T_2377; // @[AxiLoadQueue.scala 96:34:@5652.6]
  wire  _T_2379; // @[AxiLoadQueue.scala 101:36:@5660.8]
  wire  _T_2380; // @[AxiLoadQueue.scala 101:86:@5661.8]
  wire  _T_2381; // @[AxiLoadQueue.scala 101:61:@5662.8]
  wire  _T_2384; // @[AxiLoadQueue.scala 103:69:@5668.10]
  wire  _T_2385; // @[AxiLoadQueue.scala 104:31:@5669.10]
  wire  _T_2386; // @[AxiLoadQueue.scala 103:94:@5670.10]
  wire  _T_2388; // @[AxiLoadQueue.scala 103:54:@5671.10]
  wire  _T_2389; // @[AxiLoadQueue.scala 103:51:@5672.10]
  wire  _GEN_660; // @[AxiLoadQueue.scala 104:53:@5673.10]
  wire  _GEN_661; // @[AxiLoadQueue.scala 101:102:@5663.8]
  wire  _GEN_662; // @[AxiLoadQueue.scala 99:27:@5656.6]
  wire  _GEN_663; // @[AxiLoadQueue.scala 95:34:@5641.4]
  wire [4:0] _T_2402; // @[util.scala 10:8:@5684.6]
  wire [4:0] _GEN_54; // @[util.scala 10:14:@5685.6]
  wire [4:0] _T_2403; // @[util.scala 10:14:@5685.6]
  wire  _T_2404; // @[AxiLoadQueue.scala 97:56:@5686.6]
  wire  _T_2405; // @[AxiLoadQueue.scala 96:50:@5687.6]
  wire  _T_2407; // @[AxiLoadQueue.scala 96:34:@5688.6]
  wire  _T_2409; // @[AxiLoadQueue.scala 101:36:@5696.8]
  wire  _T_2410; // @[AxiLoadQueue.scala 101:86:@5697.8]
  wire  _T_2411; // @[AxiLoadQueue.scala 101:61:@5698.8]
  wire  _T_2414; // @[AxiLoadQueue.scala 103:69:@5704.10]
  wire  _T_2415; // @[AxiLoadQueue.scala 104:31:@5705.10]
  wire  _T_2416; // @[AxiLoadQueue.scala 103:94:@5706.10]
  wire  _T_2418; // @[AxiLoadQueue.scala 103:54:@5707.10]
  wire  _T_2419; // @[AxiLoadQueue.scala 103:51:@5708.10]
  wire  _GEN_680; // @[AxiLoadQueue.scala 104:53:@5709.10]
  wire  _GEN_681; // @[AxiLoadQueue.scala 101:102:@5699.8]
  wire  _GEN_682; // @[AxiLoadQueue.scala 99:27:@5692.6]
  wire  _GEN_683; // @[AxiLoadQueue.scala 95:34:@5677.4]
  wire [4:0] _T_2432; // @[util.scala 10:8:@5720.6]
  wire [4:0] _GEN_55; // @[util.scala 10:14:@5721.6]
  wire [4:0] _T_2433; // @[util.scala 10:14:@5721.6]
  wire  _T_2434; // @[AxiLoadQueue.scala 97:56:@5722.6]
  wire  _T_2435; // @[AxiLoadQueue.scala 96:50:@5723.6]
  wire  _T_2437; // @[AxiLoadQueue.scala 96:34:@5724.6]
  wire  _T_2439; // @[AxiLoadQueue.scala 101:36:@5732.8]
  wire  _T_2440; // @[AxiLoadQueue.scala 101:86:@5733.8]
  wire  _T_2441; // @[AxiLoadQueue.scala 101:61:@5734.8]
  wire  _T_2444; // @[AxiLoadQueue.scala 103:69:@5740.10]
  wire  _T_2445; // @[AxiLoadQueue.scala 104:31:@5741.10]
  wire  _T_2446; // @[AxiLoadQueue.scala 103:94:@5742.10]
  wire  _T_2448; // @[AxiLoadQueue.scala 103:54:@5743.10]
  wire  _T_2449; // @[AxiLoadQueue.scala 103:51:@5744.10]
  wire  _GEN_700; // @[AxiLoadQueue.scala 104:53:@5745.10]
  wire  _GEN_701; // @[AxiLoadQueue.scala 101:102:@5735.8]
  wire  _GEN_702; // @[AxiLoadQueue.scala 99:27:@5728.6]
  wire  _GEN_703; // @[AxiLoadQueue.scala 95:34:@5713.4]
  wire [4:0] _T_2462; // @[util.scala 10:8:@5756.6]
  wire [4:0] _GEN_56; // @[util.scala 10:14:@5757.6]
  wire [4:0] _T_2463; // @[util.scala 10:14:@5757.6]
  wire  _T_2464; // @[AxiLoadQueue.scala 97:56:@5758.6]
  wire  _T_2465; // @[AxiLoadQueue.scala 96:50:@5759.6]
  wire  _T_2467; // @[AxiLoadQueue.scala 96:34:@5760.6]
  wire  _T_2469; // @[AxiLoadQueue.scala 101:36:@5768.8]
  wire  _T_2470; // @[AxiLoadQueue.scala 101:86:@5769.8]
  wire  _T_2471; // @[AxiLoadQueue.scala 101:61:@5770.8]
  wire  _T_2474; // @[AxiLoadQueue.scala 103:69:@5776.10]
  wire  _T_2475; // @[AxiLoadQueue.scala 104:31:@5777.10]
  wire  _T_2476; // @[AxiLoadQueue.scala 103:94:@5778.10]
  wire  _T_2478; // @[AxiLoadQueue.scala 103:54:@5779.10]
  wire  _T_2479; // @[AxiLoadQueue.scala 103:51:@5780.10]
  wire  _GEN_720; // @[AxiLoadQueue.scala 104:53:@5781.10]
  wire  _GEN_721; // @[AxiLoadQueue.scala 101:102:@5771.8]
  wire  _GEN_722; // @[AxiLoadQueue.scala 99:27:@5764.6]
  wire  _GEN_723; // @[AxiLoadQueue.scala 95:34:@5749.4]
  wire [4:0] _T_2492; // @[util.scala 10:8:@5792.6]
  wire [4:0] _GEN_57; // @[util.scala 10:14:@5793.6]
  wire [4:0] _T_2493; // @[util.scala 10:14:@5793.6]
  wire  _T_2494; // @[AxiLoadQueue.scala 97:56:@5794.6]
  wire  _T_2495; // @[AxiLoadQueue.scala 96:50:@5795.6]
  wire  _T_2497; // @[AxiLoadQueue.scala 96:34:@5796.6]
  wire  _T_2499; // @[AxiLoadQueue.scala 101:36:@5804.8]
  wire  _T_2500; // @[AxiLoadQueue.scala 101:86:@5805.8]
  wire  _T_2501; // @[AxiLoadQueue.scala 101:61:@5806.8]
  wire  _T_2504; // @[AxiLoadQueue.scala 103:69:@5812.10]
  wire  _T_2505; // @[AxiLoadQueue.scala 104:31:@5813.10]
  wire  _T_2506; // @[AxiLoadQueue.scala 103:94:@5814.10]
  wire  _T_2508; // @[AxiLoadQueue.scala 103:54:@5815.10]
  wire  _T_2509; // @[AxiLoadQueue.scala 103:51:@5816.10]
  wire  _GEN_740; // @[AxiLoadQueue.scala 104:53:@5817.10]
  wire  _GEN_741; // @[AxiLoadQueue.scala 101:102:@5807.8]
  wire  _GEN_742; // @[AxiLoadQueue.scala 99:27:@5800.6]
  wire  _GEN_743; // @[AxiLoadQueue.scala 95:34:@5785.4]
  wire [4:0] _T_2522; // @[util.scala 10:8:@5828.6]
  wire [4:0] _GEN_58; // @[util.scala 10:14:@5829.6]
  wire [4:0] _T_2523; // @[util.scala 10:14:@5829.6]
  wire  _T_2524; // @[AxiLoadQueue.scala 97:56:@5830.6]
  wire  _T_2525; // @[AxiLoadQueue.scala 96:50:@5831.6]
  wire  _T_2527; // @[AxiLoadQueue.scala 96:34:@5832.6]
  wire  _T_2529; // @[AxiLoadQueue.scala 101:36:@5840.8]
  wire  _T_2530; // @[AxiLoadQueue.scala 101:86:@5841.8]
  wire  _T_2531; // @[AxiLoadQueue.scala 101:61:@5842.8]
  wire  _T_2534; // @[AxiLoadQueue.scala 103:69:@5848.10]
  wire  _T_2535; // @[AxiLoadQueue.scala 104:31:@5849.10]
  wire  _T_2536; // @[AxiLoadQueue.scala 103:94:@5850.10]
  wire  _T_2538; // @[AxiLoadQueue.scala 103:54:@5851.10]
  wire  _T_2539; // @[AxiLoadQueue.scala 103:51:@5852.10]
  wire  _GEN_760; // @[AxiLoadQueue.scala 104:53:@5853.10]
  wire  _GEN_761; // @[AxiLoadQueue.scala 101:102:@5843.8]
  wire  _GEN_762; // @[AxiLoadQueue.scala 99:27:@5836.6]
  wire  _GEN_763; // @[AxiLoadQueue.scala 95:34:@5821.4]
  wire [4:0] _T_2552; // @[util.scala 10:8:@5864.6]
  wire [4:0] _GEN_59; // @[util.scala 10:14:@5865.6]
  wire [4:0] _T_2553; // @[util.scala 10:14:@5865.6]
  wire  _T_2554; // @[AxiLoadQueue.scala 97:56:@5866.6]
  wire  _T_2555; // @[AxiLoadQueue.scala 96:50:@5867.6]
  wire  _T_2557; // @[AxiLoadQueue.scala 96:34:@5868.6]
  wire  _T_2559; // @[AxiLoadQueue.scala 101:36:@5876.8]
  wire  _T_2560; // @[AxiLoadQueue.scala 101:86:@5877.8]
  wire  _T_2561; // @[AxiLoadQueue.scala 101:61:@5878.8]
  wire  _T_2564; // @[AxiLoadQueue.scala 103:69:@5884.10]
  wire  _T_2565; // @[AxiLoadQueue.scala 104:31:@5885.10]
  wire  _T_2566; // @[AxiLoadQueue.scala 103:94:@5886.10]
  wire  _T_2568; // @[AxiLoadQueue.scala 103:54:@5887.10]
  wire  _T_2569; // @[AxiLoadQueue.scala 103:51:@5888.10]
  wire  _GEN_780; // @[AxiLoadQueue.scala 104:53:@5889.10]
  wire  _GEN_781; // @[AxiLoadQueue.scala 101:102:@5879.8]
  wire  _GEN_782; // @[AxiLoadQueue.scala 99:27:@5872.6]
  wire  _GEN_783; // @[AxiLoadQueue.scala 95:34:@5857.4]
  wire [4:0] _T_2582; // @[util.scala 10:8:@5900.6]
  wire [4:0] _GEN_60; // @[util.scala 10:14:@5901.6]
  wire [4:0] _T_2583; // @[util.scala 10:14:@5901.6]
  wire  _T_2584; // @[AxiLoadQueue.scala 97:56:@5902.6]
  wire  _T_2585; // @[AxiLoadQueue.scala 96:50:@5903.6]
  wire  _T_2587; // @[AxiLoadQueue.scala 96:34:@5904.6]
  wire  _T_2589; // @[AxiLoadQueue.scala 101:36:@5912.8]
  wire  _T_2590; // @[AxiLoadQueue.scala 101:86:@5913.8]
  wire  _T_2591; // @[AxiLoadQueue.scala 101:61:@5914.8]
  wire  _T_2594; // @[AxiLoadQueue.scala 103:69:@5920.10]
  wire  _T_2595; // @[AxiLoadQueue.scala 104:31:@5921.10]
  wire  _T_2596; // @[AxiLoadQueue.scala 103:94:@5922.10]
  wire  _T_2598; // @[AxiLoadQueue.scala 103:54:@5923.10]
  wire  _T_2599; // @[AxiLoadQueue.scala 103:51:@5924.10]
  wire  _GEN_800; // @[AxiLoadQueue.scala 104:53:@5925.10]
  wire  _GEN_801; // @[AxiLoadQueue.scala 101:102:@5915.8]
  wire  _GEN_802; // @[AxiLoadQueue.scala 99:27:@5908.6]
  wire  _GEN_803; // @[AxiLoadQueue.scala 95:34:@5893.4]
  wire [4:0] _T_2612; // @[util.scala 10:8:@5936.6]
  wire [4:0] _GEN_61; // @[util.scala 10:14:@5937.6]
  wire [4:0] _T_2613; // @[util.scala 10:14:@5937.6]
  wire  _T_2614; // @[AxiLoadQueue.scala 97:56:@5938.6]
  wire  _T_2615; // @[AxiLoadQueue.scala 96:50:@5939.6]
  wire  _T_2617; // @[AxiLoadQueue.scala 96:34:@5940.6]
  wire  _T_2619; // @[AxiLoadQueue.scala 101:36:@5948.8]
  wire  _T_2620; // @[AxiLoadQueue.scala 101:86:@5949.8]
  wire  _T_2621; // @[AxiLoadQueue.scala 101:61:@5950.8]
  wire  _T_2624; // @[AxiLoadQueue.scala 103:69:@5956.10]
  wire  _T_2625; // @[AxiLoadQueue.scala 104:31:@5957.10]
  wire  _T_2626; // @[AxiLoadQueue.scala 103:94:@5958.10]
  wire  _T_2628; // @[AxiLoadQueue.scala 103:54:@5959.10]
  wire  _T_2629; // @[AxiLoadQueue.scala 103:51:@5960.10]
  wire  _GEN_820; // @[AxiLoadQueue.scala 104:53:@5961.10]
  wire  _GEN_821; // @[AxiLoadQueue.scala 101:102:@5951.8]
  wire  _GEN_822; // @[AxiLoadQueue.scala 99:27:@5944.6]
  wire  _GEN_823; // @[AxiLoadQueue.scala 95:34:@5929.4]
  wire [4:0] _T_2642; // @[util.scala 10:8:@5972.6]
  wire [4:0] _GEN_62; // @[util.scala 10:14:@5973.6]
  wire [4:0] _T_2643; // @[util.scala 10:14:@5973.6]
  wire  _T_2644; // @[AxiLoadQueue.scala 97:56:@5974.6]
  wire  _T_2645; // @[AxiLoadQueue.scala 96:50:@5975.6]
  wire  _T_2647; // @[AxiLoadQueue.scala 96:34:@5976.6]
  wire  _T_2649; // @[AxiLoadQueue.scala 101:36:@5984.8]
  wire  _T_2650; // @[AxiLoadQueue.scala 101:86:@5985.8]
  wire  _T_2651; // @[AxiLoadQueue.scala 101:61:@5986.8]
  wire  _T_2654; // @[AxiLoadQueue.scala 103:69:@5992.10]
  wire  _T_2655; // @[AxiLoadQueue.scala 104:31:@5993.10]
  wire  _T_2656; // @[AxiLoadQueue.scala 103:94:@5994.10]
  wire  _T_2658; // @[AxiLoadQueue.scala 103:54:@5995.10]
  wire  _T_2659; // @[AxiLoadQueue.scala 103:51:@5996.10]
  wire  _GEN_840; // @[AxiLoadQueue.scala 104:53:@5997.10]
  wire  _GEN_841; // @[AxiLoadQueue.scala 101:102:@5987.8]
  wire  _GEN_842; // @[AxiLoadQueue.scala 99:27:@5980.6]
  wire  _GEN_843; // @[AxiLoadQueue.scala 95:34:@5965.4]
  wire [4:0] _T_2672; // @[util.scala 10:8:@6008.6]
  wire [4:0] _GEN_63; // @[util.scala 10:14:@6009.6]
  wire [4:0] _T_2673; // @[util.scala 10:14:@6009.6]
  wire  _T_2674; // @[AxiLoadQueue.scala 97:56:@6010.6]
  wire  _T_2675; // @[AxiLoadQueue.scala 96:50:@6011.6]
  wire  _T_2677; // @[AxiLoadQueue.scala 96:34:@6012.6]
  wire  _T_2679; // @[AxiLoadQueue.scala 101:36:@6020.8]
  wire  _T_2680; // @[AxiLoadQueue.scala 101:86:@6021.8]
  wire  _T_2681; // @[AxiLoadQueue.scala 101:61:@6022.8]
  wire  _T_2684; // @[AxiLoadQueue.scala 103:69:@6028.10]
  wire  _T_2685; // @[AxiLoadQueue.scala 104:31:@6029.10]
  wire  _T_2686; // @[AxiLoadQueue.scala 103:94:@6030.10]
  wire  _T_2688; // @[AxiLoadQueue.scala 103:54:@6031.10]
  wire  _T_2689; // @[AxiLoadQueue.scala 103:51:@6032.10]
  wire  _GEN_860; // @[AxiLoadQueue.scala 104:53:@6033.10]
  wire  _GEN_861; // @[AxiLoadQueue.scala 101:102:@6023.8]
  wire  _GEN_862; // @[AxiLoadQueue.scala 99:27:@6016.6]
  wire  _GEN_863; // @[AxiLoadQueue.scala 95:34:@6001.4]
  wire [15:0] _T_2693; // @[OneHot.scala 52:12:@6038.4]
  wire  _T_2695; // @[util.scala 60:60:@6040.4]
  wire  _T_2696; // @[util.scala 60:60:@6041.4]
  wire  _T_2697; // @[util.scala 60:60:@6042.4]
  wire  _T_2698; // @[util.scala 60:60:@6043.4]
  wire  _T_2699; // @[util.scala 60:60:@6044.4]
  wire  _T_2700; // @[util.scala 60:60:@6045.4]
  wire  _T_2701; // @[util.scala 60:60:@6046.4]
  wire  _T_2702; // @[util.scala 60:60:@6047.4]
  wire  _T_2703; // @[util.scala 60:60:@6048.4]
  wire  _T_2704; // @[util.scala 60:60:@6049.4]
  wire  _T_2705; // @[util.scala 60:60:@6050.4]
  wire  _T_2706; // @[util.scala 60:60:@6051.4]
  wire  _T_2707; // @[util.scala 60:60:@6052.4]
  wire  _T_2708; // @[util.scala 60:60:@6053.4]
  wire  _T_2709; // @[util.scala 60:60:@6054.4]
  wire  _T_2710; // @[util.scala 60:60:@6055.4]
  wire [255:0] _T_4841; // @[Mux.scala 19:72:@7579.4]
  wire [255:0] _T_4848; // @[Mux.scala 19:72:@7586.4]
  wire [511:0] _T_4849; // @[Mux.scala 19:72:@7587.4]
  wire [511:0] _T_4851; // @[Mux.scala 19:72:@7588.4]
  wire [255:0] _T_4858; // @[Mux.scala 19:72:@7595.4]
  wire [255:0] _T_4865; // @[Mux.scala 19:72:@7602.4]
  wire [511:0] _T_4866; // @[Mux.scala 19:72:@7603.4]
  wire [511:0] _T_4868; // @[Mux.scala 19:72:@7604.4]
  wire [255:0] _T_4875; // @[Mux.scala 19:72:@7611.4]
  wire [255:0] _T_4882; // @[Mux.scala 19:72:@7618.4]
  wire [511:0] _T_4883; // @[Mux.scala 19:72:@7619.4]
  wire [511:0] _T_4885; // @[Mux.scala 19:72:@7620.4]
  wire [255:0] _T_4892; // @[Mux.scala 19:72:@7627.4]
  wire [255:0] _T_4899; // @[Mux.scala 19:72:@7634.4]
  wire [511:0] _T_4900; // @[Mux.scala 19:72:@7635.4]
  wire [511:0] _T_4902; // @[Mux.scala 19:72:@7636.4]
  wire [255:0] _T_4909; // @[Mux.scala 19:72:@7643.4]
  wire [255:0] _T_4916; // @[Mux.scala 19:72:@7650.4]
  wire [511:0] _T_4917; // @[Mux.scala 19:72:@7651.4]
  wire [511:0] _T_4919; // @[Mux.scala 19:72:@7652.4]
  wire [255:0] _T_4926; // @[Mux.scala 19:72:@7659.4]
  wire [255:0] _T_4933; // @[Mux.scala 19:72:@7666.4]
  wire [511:0] _T_4934; // @[Mux.scala 19:72:@7667.4]
  wire [511:0] _T_4936; // @[Mux.scala 19:72:@7668.4]
  wire [255:0] _T_4943; // @[Mux.scala 19:72:@7675.4]
  wire [255:0] _T_4950; // @[Mux.scala 19:72:@7682.4]
  wire [511:0] _T_4951; // @[Mux.scala 19:72:@7683.4]
  wire [511:0] _T_4953; // @[Mux.scala 19:72:@7684.4]
  wire [255:0] _T_4960; // @[Mux.scala 19:72:@7691.4]
  wire [255:0] _T_4967; // @[Mux.scala 19:72:@7698.4]
  wire [511:0] _T_4968; // @[Mux.scala 19:72:@7699.4]
  wire [511:0] _T_4970; // @[Mux.scala 19:72:@7700.4]
  wire [511:0] _T_4985; // @[Mux.scala 19:72:@7715.4]
  wire [511:0] _T_4987; // @[Mux.scala 19:72:@7716.4]
  wire [511:0] _T_5002; // @[Mux.scala 19:72:@7731.4]
  wire [511:0] _T_5004; // @[Mux.scala 19:72:@7732.4]
  wire [511:0] _T_5019; // @[Mux.scala 19:72:@7747.4]
  wire [511:0] _T_5021; // @[Mux.scala 19:72:@7748.4]
  wire [511:0] _T_5036; // @[Mux.scala 19:72:@7763.4]
  wire [511:0] _T_5038; // @[Mux.scala 19:72:@7764.4]
  wire [511:0] _T_5053; // @[Mux.scala 19:72:@7779.4]
  wire [511:0] _T_5055; // @[Mux.scala 19:72:@7780.4]
  wire [511:0] _T_5070; // @[Mux.scala 19:72:@7795.4]
  wire [511:0] _T_5072; // @[Mux.scala 19:72:@7796.4]
  wire [511:0] _T_5087; // @[Mux.scala 19:72:@7811.4]
  wire [511:0] _T_5089; // @[Mux.scala 19:72:@7812.4]
  wire [511:0] _T_5104; // @[Mux.scala 19:72:@7827.4]
  wire [511:0] _T_5106; // @[Mux.scala 19:72:@7828.4]
  wire [511:0] _T_5107; // @[Mux.scala 19:72:@7829.4]
  wire [511:0] _T_5108; // @[Mux.scala 19:72:@7830.4]
  wire [511:0] _T_5109; // @[Mux.scala 19:72:@7831.4]
  wire [511:0] _T_5110; // @[Mux.scala 19:72:@7832.4]
  wire [511:0] _T_5111; // @[Mux.scala 19:72:@7833.4]
  wire [511:0] _T_5112; // @[Mux.scala 19:72:@7834.4]
  wire [511:0] _T_5113; // @[Mux.scala 19:72:@7835.4]
  wire [511:0] _T_5114; // @[Mux.scala 19:72:@7836.4]
  wire [511:0] _T_5115; // @[Mux.scala 19:72:@7837.4]
  wire [511:0] _T_5116; // @[Mux.scala 19:72:@7838.4]
  wire [511:0] _T_5117; // @[Mux.scala 19:72:@7839.4]
  wire [511:0] _T_5118; // @[Mux.scala 19:72:@7840.4]
  wire [511:0] _T_5119; // @[Mux.scala 19:72:@7841.4]
  wire [511:0] _T_5120; // @[Mux.scala 19:72:@7842.4]
  wire [511:0] _T_5121; // @[Mux.scala 19:72:@7843.4]
  wire [7:0] _T_5698; // @[Mux.scala 19:72:@8193.4]
  wire [7:0] _T_5705; // @[Mux.scala 19:72:@8200.4]
  wire [15:0] _T_5706; // @[Mux.scala 19:72:@8201.4]
  wire [15:0] _T_5708; // @[Mux.scala 19:72:@8202.4]
  wire [7:0] _T_5715; // @[Mux.scala 19:72:@8209.4]
  wire [7:0] _T_5722; // @[Mux.scala 19:72:@8216.4]
  wire [15:0] _T_5723; // @[Mux.scala 19:72:@8217.4]
  wire [15:0] _T_5725; // @[Mux.scala 19:72:@8218.4]
  wire [7:0] _T_5732; // @[Mux.scala 19:72:@8225.4]
  wire [7:0] _T_5739; // @[Mux.scala 19:72:@8232.4]
  wire [15:0] _T_5740; // @[Mux.scala 19:72:@8233.4]
  wire [15:0] _T_5742; // @[Mux.scala 19:72:@8234.4]
  wire [7:0] _T_5749; // @[Mux.scala 19:72:@8241.4]
  wire [7:0] _T_5756; // @[Mux.scala 19:72:@8248.4]
  wire [15:0] _T_5757; // @[Mux.scala 19:72:@8249.4]
  wire [15:0] _T_5759; // @[Mux.scala 19:72:@8250.4]
  wire [7:0] _T_5766; // @[Mux.scala 19:72:@8257.4]
  wire [7:0] _T_5773; // @[Mux.scala 19:72:@8264.4]
  wire [15:0] _T_5774; // @[Mux.scala 19:72:@8265.4]
  wire [15:0] _T_5776; // @[Mux.scala 19:72:@8266.4]
  wire [7:0] _T_5783; // @[Mux.scala 19:72:@8273.4]
  wire [7:0] _T_5790; // @[Mux.scala 19:72:@8280.4]
  wire [15:0] _T_5791; // @[Mux.scala 19:72:@8281.4]
  wire [15:0] _T_5793; // @[Mux.scala 19:72:@8282.4]
  wire [7:0] _T_5800; // @[Mux.scala 19:72:@8289.4]
  wire [7:0] _T_5807; // @[Mux.scala 19:72:@8296.4]
  wire [15:0] _T_5808; // @[Mux.scala 19:72:@8297.4]
  wire [15:0] _T_5810; // @[Mux.scala 19:72:@8298.4]
  wire [7:0] _T_5817; // @[Mux.scala 19:72:@8305.4]
  wire [7:0] _T_5824; // @[Mux.scala 19:72:@8312.4]
  wire [15:0] _T_5825; // @[Mux.scala 19:72:@8313.4]
  wire [15:0] _T_5827; // @[Mux.scala 19:72:@8314.4]
  wire [15:0] _T_5842; // @[Mux.scala 19:72:@8329.4]
  wire [15:0] _T_5844; // @[Mux.scala 19:72:@8330.4]
  wire [15:0] _T_5859; // @[Mux.scala 19:72:@8345.4]
  wire [15:0] _T_5861; // @[Mux.scala 19:72:@8346.4]
  wire [15:0] _T_5876; // @[Mux.scala 19:72:@8361.4]
  wire [15:0] _T_5878; // @[Mux.scala 19:72:@8362.4]
  wire [15:0] _T_5893; // @[Mux.scala 19:72:@8377.4]
  wire [15:0] _T_5895; // @[Mux.scala 19:72:@8378.4]
  wire [15:0] _T_5910; // @[Mux.scala 19:72:@8393.4]
  wire [15:0] _T_5912; // @[Mux.scala 19:72:@8394.4]
  wire [15:0] _T_5927; // @[Mux.scala 19:72:@8409.4]
  wire [15:0] _T_5929; // @[Mux.scala 19:72:@8410.4]
  wire [15:0] _T_5944; // @[Mux.scala 19:72:@8425.4]
  wire [15:0] _T_5946; // @[Mux.scala 19:72:@8426.4]
  wire [15:0] _T_5961; // @[Mux.scala 19:72:@8441.4]
  wire [15:0] _T_5963; // @[Mux.scala 19:72:@8442.4]
  wire [15:0] _T_5964; // @[Mux.scala 19:72:@8443.4]
  wire [15:0] _T_5965; // @[Mux.scala 19:72:@8444.4]
  wire [15:0] _T_5966; // @[Mux.scala 19:72:@8445.4]
  wire [15:0] _T_5967; // @[Mux.scala 19:72:@8446.4]
  wire [15:0] _T_5968; // @[Mux.scala 19:72:@8447.4]
  wire [15:0] _T_5969; // @[Mux.scala 19:72:@8448.4]
  wire [15:0] _T_5970; // @[Mux.scala 19:72:@8449.4]
  wire [15:0] _T_5971; // @[Mux.scala 19:72:@8450.4]
  wire [15:0] _T_5972; // @[Mux.scala 19:72:@8451.4]
  wire [15:0] _T_5973; // @[Mux.scala 19:72:@8452.4]
  wire [15:0] _T_5974; // @[Mux.scala 19:72:@8453.4]
  wire [15:0] _T_5975; // @[Mux.scala 19:72:@8454.4]
  wire [15:0] _T_5976; // @[Mux.scala 19:72:@8455.4]
  wire [15:0] _T_5977; // @[Mux.scala 19:72:@8456.4]
  wire [15:0] _T_5978; // @[Mux.scala 19:72:@8457.4]
  wire  _T_6119; // @[AxiLoadQueue.scala 121:105:@8493.4]
  wire  _T_6121; // @[AxiLoadQueue.scala 122:18:@8494.4]
  wire  _T_6123; // @[AxiLoadQueue.scala 122:36:@8495.4]
  wire  _T_6124; // @[AxiLoadQueue.scala 122:27:@8496.4]
  wire  _T_6126; // @[AxiLoadQueue.scala 122:52:@8497.4]
  wire  _T_6128; // @[AxiLoadQueue.scala 122:85:@8498.4]
  wire  _T_6130; // @[AxiLoadQueue.scala 122:103:@8499.4]
  wire  _T_6131; // @[AxiLoadQueue.scala 122:94:@8500.4]
  wire  _T_6133; // @[AxiLoadQueue.scala 122:70:@8501.4]
  wire  _T_6134; // @[AxiLoadQueue.scala 122:67:@8502.4]
  wire  validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 121:91:@8503.4]
  wire  _T_6138; // @[AxiLoadQueue.scala 122:18:@8505.4]
  wire  _T_6140; // @[AxiLoadQueue.scala 122:36:@8506.4]
  wire  _T_6141; // @[AxiLoadQueue.scala 122:27:@8507.4]
  wire  _T_6145; // @[AxiLoadQueue.scala 122:85:@8509.4]
  wire  _T_6147; // @[AxiLoadQueue.scala 122:103:@8510.4]
  wire  _T_6148; // @[AxiLoadQueue.scala 122:94:@8511.4]
  wire  _T_6150; // @[AxiLoadQueue.scala 122:70:@8512.4]
  wire  _T_6151; // @[AxiLoadQueue.scala 122:67:@8513.4]
  wire  validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 121:91:@8514.4]
  wire  _T_6155; // @[AxiLoadQueue.scala 122:18:@8516.4]
  wire  _T_6157; // @[AxiLoadQueue.scala 122:36:@8517.4]
  wire  _T_6158; // @[AxiLoadQueue.scala 122:27:@8518.4]
  wire  _T_6162; // @[AxiLoadQueue.scala 122:85:@8520.4]
  wire  _T_6164; // @[AxiLoadQueue.scala 122:103:@8521.4]
  wire  _T_6165; // @[AxiLoadQueue.scala 122:94:@8522.4]
  wire  _T_6167; // @[AxiLoadQueue.scala 122:70:@8523.4]
  wire  _T_6168; // @[AxiLoadQueue.scala 122:67:@8524.4]
  wire  validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 121:91:@8525.4]
  wire  _T_6172; // @[AxiLoadQueue.scala 122:18:@8527.4]
  wire  _T_6174; // @[AxiLoadQueue.scala 122:36:@8528.4]
  wire  _T_6175; // @[AxiLoadQueue.scala 122:27:@8529.4]
  wire  _T_6179; // @[AxiLoadQueue.scala 122:85:@8531.4]
  wire  _T_6181; // @[AxiLoadQueue.scala 122:103:@8532.4]
  wire  _T_6182; // @[AxiLoadQueue.scala 122:94:@8533.4]
  wire  _T_6184; // @[AxiLoadQueue.scala 122:70:@8534.4]
  wire  _T_6185; // @[AxiLoadQueue.scala 122:67:@8535.4]
  wire  validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 121:91:@8536.4]
  wire  _T_6189; // @[AxiLoadQueue.scala 122:18:@8538.4]
  wire  _T_6191; // @[AxiLoadQueue.scala 122:36:@8539.4]
  wire  _T_6192; // @[AxiLoadQueue.scala 122:27:@8540.4]
  wire  _T_6196; // @[AxiLoadQueue.scala 122:85:@8542.4]
  wire  _T_6198; // @[AxiLoadQueue.scala 122:103:@8543.4]
  wire  _T_6199; // @[AxiLoadQueue.scala 122:94:@8544.4]
  wire  _T_6201; // @[AxiLoadQueue.scala 122:70:@8545.4]
  wire  _T_6202; // @[AxiLoadQueue.scala 122:67:@8546.4]
  wire  validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 121:91:@8547.4]
  wire  _T_6206; // @[AxiLoadQueue.scala 122:18:@8549.4]
  wire  _T_6208; // @[AxiLoadQueue.scala 122:36:@8550.4]
  wire  _T_6209; // @[AxiLoadQueue.scala 122:27:@8551.4]
  wire  _T_6213; // @[AxiLoadQueue.scala 122:85:@8553.4]
  wire  _T_6215; // @[AxiLoadQueue.scala 122:103:@8554.4]
  wire  _T_6216; // @[AxiLoadQueue.scala 122:94:@8555.4]
  wire  _T_6218; // @[AxiLoadQueue.scala 122:70:@8556.4]
  wire  _T_6219; // @[AxiLoadQueue.scala 122:67:@8557.4]
  wire  validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 121:91:@8558.4]
  wire  _T_6223; // @[AxiLoadQueue.scala 122:18:@8560.4]
  wire  _T_6225; // @[AxiLoadQueue.scala 122:36:@8561.4]
  wire  _T_6226; // @[AxiLoadQueue.scala 122:27:@8562.4]
  wire  _T_6230; // @[AxiLoadQueue.scala 122:85:@8564.4]
  wire  _T_6232; // @[AxiLoadQueue.scala 122:103:@8565.4]
  wire  _T_6233; // @[AxiLoadQueue.scala 122:94:@8566.4]
  wire  _T_6235; // @[AxiLoadQueue.scala 122:70:@8567.4]
  wire  _T_6236; // @[AxiLoadQueue.scala 122:67:@8568.4]
  wire  validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 121:91:@8569.4]
  wire  _T_6240; // @[AxiLoadQueue.scala 122:18:@8571.4]
  wire  _T_6242; // @[AxiLoadQueue.scala 122:36:@8572.4]
  wire  _T_6243; // @[AxiLoadQueue.scala 122:27:@8573.4]
  wire  _T_6247; // @[AxiLoadQueue.scala 122:85:@8575.4]
  wire  _T_6249; // @[AxiLoadQueue.scala 122:103:@8576.4]
  wire  _T_6250; // @[AxiLoadQueue.scala 122:94:@8577.4]
  wire  _T_6252; // @[AxiLoadQueue.scala 122:70:@8578.4]
  wire  _T_6253; // @[AxiLoadQueue.scala 122:67:@8579.4]
  wire  validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 121:91:@8580.4]
  wire  _T_6257; // @[AxiLoadQueue.scala 122:18:@8582.4]
  wire  _T_6259; // @[AxiLoadQueue.scala 122:36:@8583.4]
  wire  _T_6260; // @[AxiLoadQueue.scala 122:27:@8584.4]
  wire  _T_6264; // @[AxiLoadQueue.scala 122:85:@8586.4]
  wire  _T_6266; // @[AxiLoadQueue.scala 122:103:@8587.4]
  wire  _T_6267; // @[AxiLoadQueue.scala 122:94:@8588.4]
  wire  _T_6269; // @[AxiLoadQueue.scala 122:70:@8589.4]
  wire  _T_6270; // @[AxiLoadQueue.scala 122:67:@8590.4]
  wire  validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 121:91:@8591.4]
  wire  _T_6274; // @[AxiLoadQueue.scala 122:18:@8593.4]
  wire  _T_6276; // @[AxiLoadQueue.scala 122:36:@8594.4]
  wire  _T_6277; // @[AxiLoadQueue.scala 122:27:@8595.4]
  wire  _T_6281; // @[AxiLoadQueue.scala 122:85:@8597.4]
  wire  _T_6283; // @[AxiLoadQueue.scala 122:103:@8598.4]
  wire  _T_6284; // @[AxiLoadQueue.scala 122:94:@8599.4]
  wire  _T_6286; // @[AxiLoadQueue.scala 122:70:@8600.4]
  wire  _T_6287; // @[AxiLoadQueue.scala 122:67:@8601.4]
  wire  validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 121:91:@8602.4]
  wire  _T_6291; // @[AxiLoadQueue.scala 122:18:@8604.4]
  wire  _T_6293; // @[AxiLoadQueue.scala 122:36:@8605.4]
  wire  _T_6294; // @[AxiLoadQueue.scala 122:27:@8606.4]
  wire  _T_6298; // @[AxiLoadQueue.scala 122:85:@8608.4]
  wire  _T_6300; // @[AxiLoadQueue.scala 122:103:@8609.4]
  wire  _T_6301; // @[AxiLoadQueue.scala 122:94:@8610.4]
  wire  _T_6303; // @[AxiLoadQueue.scala 122:70:@8611.4]
  wire  _T_6304; // @[AxiLoadQueue.scala 122:67:@8612.4]
  wire  validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 121:91:@8613.4]
  wire  _T_6308; // @[AxiLoadQueue.scala 122:18:@8615.4]
  wire  _T_6310; // @[AxiLoadQueue.scala 122:36:@8616.4]
  wire  _T_6311; // @[AxiLoadQueue.scala 122:27:@8617.4]
  wire  _T_6315; // @[AxiLoadQueue.scala 122:85:@8619.4]
  wire  _T_6317; // @[AxiLoadQueue.scala 122:103:@8620.4]
  wire  _T_6318; // @[AxiLoadQueue.scala 122:94:@8621.4]
  wire  _T_6320; // @[AxiLoadQueue.scala 122:70:@8622.4]
  wire  _T_6321; // @[AxiLoadQueue.scala 122:67:@8623.4]
  wire  validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 121:91:@8624.4]
  wire  _T_6325; // @[AxiLoadQueue.scala 122:18:@8626.4]
  wire  _T_6327; // @[AxiLoadQueue.scala 122:36:@8627.4]
  wire  _T_6328; // @[AxiLoadQueue.scala 122:27:@8628.4]
  wire  _T_6332; // @[AxiLoadQueue.scala 122:85:@8630.4]
  wire  _T_6334; // @[AxiLoadQueue.scala 122:103:@8631.4]
  wire  _T_6335; // @[AxiLoadQueue.scala 122:94:@8632.4]
  wire  _T_6337; // @[AxiLoadQueue.scala 122:70:@8633.4]
  wire  _T_6338; // @[AxiLoadQueue.scala 122:67:@8634.4]
  wire  validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 121:91:@8635.4]
  wire  _T_6342; // @[AxiLoadQueue.scala 122:18:@8637.4]
  wire  _T_6344; // @[AxiLoadQueue.scala 122:36:@8638.4]
  wire  _T_6345; // @[AxiLoadQueue.scala 122:27:@8639.4]
  wire  _T_6349; // @[AxiLoadQueue.scala 122:85:@8641.4]
  wire  _T_6351; // @[AxiLoadQueue.scala 122:103:@8642.4]
  wire  _T_6352; // @[AxiLoadQueue.scala 122:94:@8643.4]
  wire  _T_6354; // @[AxiLoadQueue.scala 122:70:@8644.4]
  wire  _T_6355; // @[AxiLoadQueue.scala 122:67:@8645.4]
  wire  validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 121:91:@8646.4]
  wire  _T_6359; // @[AxiLoadQueue.scala 122:18:@8648.4]
  wire  _T_6361; // @[AxiLoadQueue.scala 122:36:@8649.4]
  wire  _T_6362; // @[AxiLoadQueue.scala 122:27:@8650.4]
  wire  _T_6366; // @[AxiLoadQueue.scala 122:85:@8652.4]
  wire  _T_6368; // @[AxiLoadQueue.scala 122:103:@8653.4]
  wire  _T_6369; // @[AxiLoadQueue.scala 122:94:@8654.4]
  wire  _T_6371; // @[AxiLoadQueue.scala 122:70:@8655.4]
  wire  _T_6372; // @[AxiLoadQueue.scala 122:67:@8656.4]
  wire  validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 121:91:@8657.4]
  wire  validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 121:91:@8668.4]
  wire  storesToCheck_0_0; // @[AxiLoadQueue.scala 130:10:@8695.4]
  wire  _T_7660; // @[AxiLoadQueue.scala 130:81:@8698.4]
  wire  _T_7661; // @[AxiLoadQueue.scala 130:72:@8699.4]
  wire  _T_7663; // @[AxiLoadQueue.scala 131:33:@8700.4]
  wire  _T_7666; // @[AxiLoadQueue.scala 131:41:@8702.4]
  wire  _T_7668; // @[AxiLoadQueue.scala 131:9:@8703.4]
  wire  storesToCheck_0_1; // @[AxiLoadQueue.scala 130:10:@8704.4]
  wire  _T_7674; // @[AxiLoadQueue.scala 130:81:@8707.4]
  wire  _T_7675; // @[AxiLoadQueue.scala 130:72:@8708.4]
  wire  _T_7677; // @[AxiLoadQueue.scala 131:33:@8709.4]
  wire  _T_7680; // @[AxiLoadQueue.scala 131:41:@8711.4]
  wire  _T_7682; // @[AxiLoadQueue.scala 131:9:@8712.4]
  wire  storesToCheck_0_2; // @[AxiLoadQueue.scala 130:10:@8713.4]
  wire  _T_7688; // @[AxiLoadQueue.scala 130:81:@8716.4]
  wire  _T_7689; // @[AxiLoadQueue.scala 130:72:@8717.4]
  wire  _T_7691; // @[AxiLoadQueue.scala 131:33:@8718.4]
  wire  _T_7694; // @[AxiLoadQueue.scala 131:41:@8720.4]
  wire  _T_7696; // @[AxiLoadQueue.scala 131:9:@8721.4]
  wire  storesToCheck_0_3; // @[AxiLoadQueue.scala 130:10:@8722.4]
  wire  _T_7702; // @[AxiLoadQueue.scala 130:81:@8725.4]
  wire  _T_7703; // @[AxiLoadQueue.scala 130:72:@8726.4]
  wire  _T_7705; // @[AxiLoadQueue.scala 131:33:@8727.4]
  wire  _T_7708; // @[AxiLoadQueue.scala 131:41:@8729.4]
  wire  _T_7710; // @[AxiLoadQueue.scala 131:9:@8730.4]
  wire  storesToCheck_0_4; // @[AxiLoadQueue.scala 130:10:@8731.4]
  wire  _T_7716; // @[AxiLoadQueue.scala 130:81:@8734.4]
  wire  _T_7717; // @[AxiLoadQueue.scala 130:72:@8735.4]
  wire  _T_7719; // @[AxiLoadQueue.scala 131:33:@8736.4]
  wire  _T_7722; // @[AxiLoadQueue.scala 131:41:@8738.4]
  wire  _T_7724; // @[AxiLoadQueue.scala 131:9:@8739.4]
  wire  storesToCheck_0_5; // @[AxiLoadQueue.scala 130:10:@8740.4]
  wire  _T_7730; // @[AxiLoadQueue.scala 130:81:@8743.4]
  wire  _T_7731; // @[AxiLoadQueue.scala 130:72:@8744.4]
  wire  _T_7733; // @[AxiLoadQueue.scala 131:33:@8745.4]
  wire  _T_7736; // @[AxiLoadQueue.scala 131:41:@8747.4]
  wire  _T_7738; // @[AxiLoadQueue.scala 131:9:@8748.4]
  wire  storesToCheck_0_6; // @[AxiLoadQueue.scala 130:10:@8749.4]
  wire  _T_7744; // @[AxiLoadQueue.scala 130:81:@8752.4]
  wire  _T_7745; // @[AxiLoadQueue.scala 130:72:@8753.4]
  wire  _T_7747; // @[AxiLoadQueue.scala 131:33:@8754.4]
  wire  _T_7750; // @[AxiLoadQueue.scala 131:41:@8756.4]
  wire  _T_7752; // @[AxiLoadQueue.scala 131:9:@8757.4]
  wire  storesToCheck_0_7; // @[AxiLoadQueue.scala 130:10:@8758.4]
  wire  _T_7758; // @[AxiLoadQueue.scala 130:81:@8761.4]
  wire  _T_7759; // @[AxiLoadQueue.scala 130:72:@8762.4]
  wire  _T_7761; // @[AxiLoadQueue.scala 131:33:@8763.4]
  wire  _T_7764; // @[AxiLoadQueue.scala 131:41:@8765.4]
  wire  _T_7766; // @[AxiLoadQueue.scala 131:9:@8766.4]
  wire  storesToCheck_0_8; // @[AxiLoadQueue.scala 130:10:@8767.4]
  wire  _T_7772; // @[AxiLoadQueue.scala 130:81:@8770.4]
  wire  _T_7773; // @[AxiLoadQueue.scala 130:72:@8771.4]
  wire  _T_7775; // @[AxiLoadQueue.scala 131:33:@8772.4]
  wire  _T_7778; // @[AxiLoadQueue.scala 131:41:@8774.4]
  wire  _T_7780; // @[AxiLoadQueue.scala 131:9:@8775.4]
  wire  storesToCheck_0_9; // @[AxiLoadQueue.scala 130:10:@8776.4]
  wire  _T_7786; // @[AxiLoadQueue.scala 130:81:@8779.4]
  wire  _T_7787; // @[AxiLoadQueue.scala 130:72:@8780.4]
  wire  _T_7789; // @[AxiLoadQueue.scala 131:33:@8781.4]
  wire  _T_7792; // @[AxiLoadQueue.scala 131:41:@8783.4]
  wire  _T_7794; // @[AxiLoadQueue.scala 131:9:@8784.4]
  wire  storesToCheck_0_10; // @[AxiLoadQueue.scala 130:10:@8785.4]
  wire  _T_7800; // @[AxiLoadQueue.scala 130:81:@8788.4]
  wire  _T_7801; // @[AxiLoadQueue.scala 130:72:@8789.4]
  wire  _T_7803; // @[AxiLoadQueue.scala 131:33:@8790.4]
  wire  _T_7806; // @[AxiLoadQueue.scala 131:41:@8792.4]
  wire  _T_7808; // @[AxiLoadQueue.scala 131:9:@8793.4]
  wire  storesToCheck_0_11; // @[AxiLoadQueue.scala 130:10:@8794.4]
  wire  _T_7814; // @[AxiLoadQueue.scala 130:81:@8797.4]
  wire  _T_7815; // @[AxiLoadQueue.scala 130:72:@8798.4]
  wire  _T_7817; // @[AxiLoadQueue.scala 131:33:@8799.4]
  wire  _T_7820; // @[AxiLoadQueue.scala 131:41:@8801.4]
  wire  _T_7822; // @[AxiLoadQueue.scala 131:9:@8802.4]
  wire  storesToCheck_0_12; // @[AxiLoadQueue.scala 130:10:@8803.4]
  wire  _T_7828; // @[AxiLoadQueue.scala 130:81:@8806.4]
  wire  _T_7829; // @[AxiLoadQueue.scala 130:72:@8807.4]
  wire  _T_7831; // @[AxiLoadQueue.scala 131:33:@8808.4]
  wire  _T_7834; // @[AxiLoadQueue.scala 131:41:@8810.4]
  wire  _T_7836; // @[AxiLoadQueue.scala 131:9:@8811.4]
  wire  storesToCheck_0_13; // @[AxiLoadQueue.scala 130:10:@8812.4]
  wire  _T_7842; // @[AxiLoadQueue.scala 130:81:@8815.4]
  wire  _T_7843; // @[AxiLoadQueue.scala 130:72:@8816.4]
  wire  _T_7845; // @[AxiLoadQueue.scala 131:33:@8817.4]
  wire  _T_7848; // @[AxiLoadQueue.scala 131:41:@8819.4]
  wire  _T_7850; // @[AxiLoadQueue.scala 131:9:@8820.4]
  wire  storesToCheck_0_14; // @[AxiLoadQueue.scala 130:10:@8821.4]
  wire  _T_7856; // @[AxiLoadQueue.scala 130:81:@8824.4]
  wire  storesToCheck_0_15; // @[AxiLoadQueue.scala 130:10:@8830.4]
  wire  storesToCheck_1_0; // @[AxiLoadQueue.scala 130:10:@8872.4]
  wire  _T_7906; // @[AxiLoadQueue.scala 130:81:@8875.4]
  wire  _T_7907; // @[AxiLoadQueue.scala 130:72:@8876.4]
  wire  _T_7909; // @[AxiLoadQueue.scala 131:33:@8877.4]
  wire  _T_7912; // @[AxiLoadQueue.scala 131:41:@8879.4]
  wire  _T_7914; // @[AxiLoadQueue.scala 131:9:@8880.4]
  wire  storesToCheck_1_1; // @[AxiLoadQueue.scala 130:10:@8881.4]
  wire  _T_7920; // @[AxiLoadQueue.scala 130:81:@8884.4]
  wire  _T_7921; // @[AxiLoadQueue.scala 130:72:@8885.4]
  wire  _T_7923; // @[AxiLoadQueue.scala 131:33:@8886.4]
  wire  _T_7926; // @[AxiLoadQueue.scala 131:41:@8888.4]
  wire  _T_7928; // @[AxiLoadQueue.scala 131:9:@8889.4]
  wire  storesToCheck_1_2; // @[AxiLoadQueue.scala 130:10:@8890.4]
  wire  _T_7934; // @[AxiLoadQueue.scala 130:81:@8893.4]
  wire  _T_7935; // @[AxiLoadQueue.scala 130:72:@8894.4]
  wire  _T_7937; // @[AxiLoadQueue.scala 131:33:@8895.4]
  wire  _T_7940; // @[AxiLoadQueue.scala 131:41:@8897.4]
  wire  _T_7942; // @[AxiLoadQueue.scala 131:9:@8898.4]
  wire  storesToCheck_1_3; // @[AxiLoadQueue.scala 130:10:@8899.4]
  wire  _T_7948; // @[AxiLoadQueue.scala 130:81:@8902.4]
  wire  _T_7949; // @[AxiLoadQueue.scala 130:72:@8903.4]
  wire  _T_7951; // @[AxiLoadQueue.scala 131:33:@8904.4]
  wire  _T_7954; // @[AxiLoadQueue.scala 131:41:@8906.4]
  wire  _T_7956; // @[AxiLoadQueue.scala 131:9:@8907.4]
  wire  storesToCheck_1_4; // @[AxiLoadQueue.scala 130:10:@8908.4]
  wire  _T_7962; // @[AxiLoadQueue.scala 130:81:@8911.4]
  wire  _T_7963; // @[AxiLoadQueue.scala 130:72:@8912.4]
  wire  _T_7965; // @[AxiLoadQueue.scala 131:33:@8913.4]
  wire  _T_7968; // @[AxiLoadQueue.scala 131:41:@8915.4]
  wire  _T_7970; // @[AxiLoadQueue.scala 131:9:@8916.4]
  wire  storesToCheck_1_5; // @[AxiLoadQueue.scala 130:10:@8917.4]
  wire  _T_7976; // @[AxiLoadQueue.scala 130:81:@8920.4]
  wire  _T_7977; // @[AxiLoadQueue.scala 130:72:@8921.4]
  wire  _T_7979; // @[AxiLoadQueue.scala 131:33:@8922.4]
  wire  _T_7982; // @[AxiLoadQueue.scala 131:41:@8924.4]
  wire  _T_7984; // @[AxiLoadQueue.scala 131:9:@8925.4]
  wire  storesToCheck_1_6; // @[AxiLoadQueue.scala 130:10:@8926.4]
  wire  _T_7990; // @[AxiLoadQueue.scala 130:81:@8929.4]
  wire  _T_7991; // @[AxiLoadQueue.scala 130:72:@8930.4]
  wire  _T_7993; // @[AxiLoadQueue.scala 131:33:@8931.4]
  wire  _T_7996; // @[AxiLoadQueue.scala 131:41:@8933.4]
  wire  _T_7998; // @[AxiLoadQueue.scala 131:9:@8934.4]
  wire  storesToCheck_1_7; // @[AxiLoadQueue.scala 130:10:@8935.4]
  wire  _T_8004; // @[AxiLoadQueue.scala 130:81:@8938.4]
  wire  _T_8005; // @[AxiLoadQueue.scala 130:72:@8939.4]
  wire  _T_8007; // @[AxiLoadQueue.scala 131:33:@8940.4]
  wire  _T_8010; // @[AxiLoadQueue.scala 131:41:@8942.4]
  wire  _T_8012; // @[AxiLoadQueue.scala 131:9:@8943.4]
  wire  storesToCheck_1_8; // @[AxiLoadQueue.scala 130:10:@8944.4]
  wire  _T_8018; // @[AxiLoadQueue.scala 130:81:@8947.4]
  wire  _T_8019; // @[AxiLoadQueue.scala 130:72:@8948.4]
  wire  _T_8021; // @[AxiLoadQueue.scala 131:33:@8949.4]
  wire  _T_8024; // @[AxiLoadQueue.scala 131:41:@8951.4]
  wire  _T_8026; // @[AxiLoadQueue.scala 131:9:@8952.4]
  wire  storesToCheck_1_9; // @[AxiLoadQueue.scala 130:10:@8953.4]
  wire  _T_8032; // @[AxiLoadQueue.scala 130:81:@8956.4]
  wire  _T_8033; // @[AxiLoadQueue.scala 130:72:@8957.4]
  wire  _T_8035; // @[AxiLoadQueue.scala 131:33:@8958.4]
  wire  _T_8038; // @[AxiLoadQueue.scala 131:41:@8960.4]
  wire  _T_8040; // @[AxiLoadQueue.scala 131:9:@8961.4]
  wire  storesToCheck_1_10; // @[AxiLoadQueue.scala 130:10:@8962.4]
  wire  _T_8046; // @[AxiLoadQueue.scala 130:81:@8965.4]
  wire  _T_8047; // @[AxiLoadQueue.scala 130:72:@8966.4]
  wire  _T_8049; // @[AxiLoadQueue.scala 131:33:@8967.4]
  wire  _T_8052; // @[AxiLoadQueue.scala 131:41:@8969.4]
  wire  _T_8054; // @[AxiLoadQueue.scala 131:9:@8970.4]
  wire  storesToCheck_1_11; // @[AxiLoadQueue.scala 130:10:@8971.4]
  wire  _T_8060; // @[AxiLoadQueue.scala 130:81:@8974.4]
  wire  _T_8061; // @[AxiLoadQueue.scala 130:72:@8975.4]
  wire  _T_8063; // @[AxiLoadQueue.scala 131:33:@8976.4]
  wire  _T_8066; // @[AxiLoadQueue.scala 131:41:@8978.4]
  wire  _T_8068; // @[AxiLoadQueue.scala 131:9:@8979.4]
  wire  storesToCheck_1_12; // @[AxiLoadQueue.scala 130:10:@8980.4]
  wire  _T_8074; // @[AxiLoadQueue.scala 130:81:@8983.4]
  wire  _T_8075; // @[AxiLoadQueue.scala 130:72:@8984.4]
  wire  _T_8077; // @[AxiLoadQueue.scala 131:33:@8985.4]
  wire  _T_8080; // @[AxiLoadQueue.scala 131:41:@8987.4]
  wire  _T_8082; // @[AxiLoadQueue.scala 131:9:@8988.4]
  wire  storesToCheck_1_13; // @[AxiLoadQueue.scala 130:10:@8989.4]
  wire  _T_8088; // @[AxiLoadQueue.scala 130:81:@8992.4]
  wire  _T_8089; // @[AxiLoadQueue.scala 130:72:@8993.4]
  wire  _T_8091; // @[AxiLoadQueue.scala 131:33:@8994.4]
  wire  _T_8094; // @[AxiLoadQueue.scala 131:41:@8996.4]
  wire  _T_8096; // @[AxiLoadQueue.scala 131:9:@8997.4]
  wire  storesToCheck_1_14; // @[AxiLoadQueue.scala 130:10:@8998.4]
  wire  _T_8102; // @[AxiLoadQueue.scala 130:81:@9001.4]
  wire  storesToCheck_1_15; // @[AxiLoadQueue.scala 130:10:@9007.4]
  wire  storesToCheck_2_0; // @[AxiLoadQueue.scala 130:10:@9049.4]
  wire  _T_8152; // @[AxiLoadQueue.scala 130:81:@9052.4]
  wire  _T_8153; // @[AxiLoadQueue.scala 130:72:@9053.4]
  wire  _T_8155; // @[AxiLoadQueue.scala 131:33:@9054.4]
  wire  _T_8158; // @[AxiLoadQueue.scala 131:41:@9056.4]
  wire  _T_8160; // @[AxiLoadQueue.scala 131:9:@9057.4]
  wire  storesToCheck_2_1; // @[AxiLoadQueue.scala 130:10:@9058.4]
  wire  _T_8166; // @[AxiLoadQueue.scala 130:81:@9061.4]
  wire  _T_8167; // @[AxiLoadQueue.scala 130:72:@9062.4]
  wire  _T_8169; // @[AxiLoadQueue.scala 131:33:@9063.4]
  wire  _T_8172; // @[AxiLoadQueue.scala 131:41:@9065.4]
  wire  _T_8174; // @[AxiLoadQueue.scala 131:9:@9066.4]
  wire  storesToCheck_2_2; // @[AxiLoadQueue.scala 130:10:@9067.4]
  wire  _T_8180; // @[AxiLoadQueue.scala 130:81:@9070.4]
  wire  _T_8181; // @[AxiLoadQueue.scala 130:72:@9071.4]
  wire  _T_8183; // @[AxiLoadQueue.scala 131:33:@9072.4]
  wire  _T_8186; // @[AxiLoadQueue.scala 131:41:@9074.4]
  wire  _T_8188; // @[AxiLoadQueue.scala 131:9:@9075.4]
  wire  storesToCheck_2_3; // @[AxiLoadQueue.scala 130:10:@9076.4]
  wire  _T_8194; // @[AxiLoadQueue.scala 130:81:@9079.4]
  wire  _T_8195; // @[AxiLoadQueue.scala 130:72:@9080.4]
  wire  _T_8197; // @[AxiLoadQueue.scala 131:33:@9081.4]
  wire  _T_8200; // @[AxiLoadQueue.scala 131:41:@9083.4]
  wire  _T_8202; // @[AxiLoadQueue.scala 131:9:@9084.4]
  wire  storesToCheck_2_4; // @[AxiLoadQueue.scala 130:10:@9085.4]
  wire  _T_8208; // @[AxiLoadQueue.scala 130:81:@9088.4]
  wire  _T_8209; // @[AxiLoadQueue.scala 130:72:@9089.4]
  wire  _T_8211; // @[AxiLoadQueue.scala 131:33:@9090.4]
  wire  _T_8214; // @[AxiLoadQueue.scala 131:41:@9092.4]
  wire  _T_8216; // @[AxiLoadQueue.scala 131:9:@9093.4]
  wire  storesToCheck_2_5; // @[AxiLoadQueue.scala 130:10:@9094.4]
  wire  _T_8222; // @[AxiLoadQueue.scala 130:81:@9097.4]
  wire  _T_8223; // @[AxiLoadQueue.scala 130:72:@9098.4]
  wire  _T_8225; // @[AxiLoadQueue.scala 131:33:@9099.4]
  wire  _T_8228; // @[AxiLoadQueue.scala 131:41:@9101.4]
  wire  _T_8230; // @[AxiLoadQueue.scala 131:9:@9102.4]
  wire  storesToCheck_2_6; // @[AxiLoadQueue.scala 130:10:@9103.4]
  wire  _T_8236; // @[AxiLoadQueue.scala 130:81:@9106.4]
  wire  _T_8237; // @[AxiLoadQueue.scala 130:72:@9107.4]
  wire  _T_8239; // @[AxiLoadQueue.scala 131:33:@9108.4]
  wire  _T_8242; // @[AxiLoadQueue.scala 131:41:@9110.4]
  wire  _T_8244; // @[AxiLoadQueue.scala 131:9:@9111.4]
  wire  storesToCheck_2_7; // @[AxiLoadQueue.scala 130:10:@9112.4]
  wire  _T_8250; // @[AxiLoadQueue.scala 130:81:@9115.4]
  wire  _T_8251; // @[AxiLoadQueue.scala 130:72:@9116.4]
  wire  _T_8253; // @[AxiLoadQueue.scala 131:33:@9117.4]
  wire  _T_8256; // @[AxiLoadQueue.scala 131:41:@9119.4]
  wire  _T_8258; // @[AxiLoadQueue.scala 131:9:@9120.4]
  wire  storesToCheck_2_8; // @[AxiLoadQueue.scala 130:10:@9121.4]
  wire  _T_8264; // @[AxiLoadQueue.scala 130:81:@9124.4]
  wire  _T_8265; // @[AxiLoadQueue.scala 130:72:@9125.4]
  wire  _T_8267; // @[AxiLoadQueue.scala 131:33:@9126.4]
  wire  _T_8270; // @[AxiLoadQueue.scala 131:41:@9128.4]
  wire  _T_8272; // @[AxiLoadQueue.scala 131:9:@9129.4]
  wire  storesToCheck_2_9; // @[AxiLoadQueue.scala 130:10:@9130.4]
  wire  _T_8278; // @[AxiLoadQueue.scala 130:81:@9133.4]
  wire  _T_8279; // @[AxiLoadQueue.scala 130:72:@9134.4]
  wire  _T_8281; // @[AxiLoadQueue.scala 131:33:@9135.4]
  wire  _T_8284; // @[AxiLoadQueue.scala 131:41:@9137.4]
  wire  _T_8286; // @[AxiLoadQueue.scala 131:9:@9138.4]
  wire  storesToCheck_2_10; // @[AxiLoadQueue.scala 130:10:@9139.4]
  wire  _T_8292; // @[AxiLoadQueue.scala 130:81:@9142.4]
  wire  _T_8293; // @[AxiLoadQueue.scala 130:72:@9143.4]
  wire  _T_8295; // @[AxiLoadQueue.scala 131:33:@9144.4]
  wire  _T_8298; // @[AxiLoadQueue.scala 131:41:@9146.4]
  wire  _T_8300; // @[AxiLoadQueue.scala 131:9:@9147.4]
  wire  storesToCheck_2_11; // @[AxiLoadQueue.scala 130:10:@9148.4]
  wire  _T_8306; // @[AxiLoadQueue.scala 130:81:@9151.4]
  wire  _T_8307; // @[AxiLoadQueue.scala 130:72:@9152.4]
  wire  _T_8309; // @[AxiLoadQueue.scala 131:33:@9153.4]
  wire  _T_8312; // @[AxiLoadQueue.scala 131:41:@9155.4]
  wire  _T_8314; // @[AxiLoadQueue.scala 131:9:@9156.4]
  wire  storesToCheck_2_12; // @[AxiLoadQueue.scala 130:10:@9157.4]
  wire  _T_8320; // @[AxiLoadQueue.scala 130:81:@9160.4]
  wire  _T_8321; // @[AxiLoadQueue.scala 130:72:@9161.4]
  wire  _T_8323; // @[AxiLoadQueue.scala 131:33:@9162.4]
  wire  _T_8326; // @[AxiLoadQueue.scala 131:41:@9164.4]
  wire  _T_8328; // @[AxiLoadQueue.scala 131:9:@9165.4]
  wire  storesToCheck_2_13; // @[AxiLoadQueue.scala 130:10:@9166.4]
  wire  _T_8334; // @[AxiLoadQueue.scala 130:81:@9169.4]
  wire  _T_8335; // @[AxiLoadQueue.scala 130:72:@9170.4]
  wire  _T_8337; // @[AxiLoadQueue.scala 131:33:@9171.4]
  wire  _T_8340; // @[AxiLoadQueue.scala 131:41:@9173.4]
  wire  _T_8342; // @[AxiLoadQueue.scala 131:9:@9174.4]
  wire  storesToCheck_2_14; // @[AxiLoadQueue.scala 130:10:@9175.4]
  wire  _T_8348; // @[AxiLoadQueue.scala 130:81:@9178.4]
  wire  storesToCheck_2_15; // @[AxiLoadQueue.scala 130:10:@9184.4]
  wire  storesToCheck_3_0; // @[AxiLoadQueue.scala 130:10:@9226.4]
  wire  _T_8398; // @[AxiLoadQueue.scala 130:81:@9229.4]
  wire  _T_8399; // @[AxiLoadQueue.scala 130:72:@9230.4]
  wire  _T_8401; // @[AxiLoadQueue.scala 131:33:@9231.4]
  wire  _T_8404; // @[AxiLoadQueue.scala 131:41:@9233.4]
  wire  _T_8406; // @[AxiLoadQueue.scala 131:9:@9234.4]
  wire  storesToCheck_3_1; // @[AxiLoadQueue.scala 130:10:@9235.4]
  wire  _T_8412; // @[AxiLoadQueue.scala 130:81:@9238.4]
  wire  _T_8413; // @[AxiLoadQueue.scala 130:72:@9239.4]
  wire  _T_8415; // @[AxiLoadQueue.scala 131:33:@9240.4]
  wire  _T_8418; // @[AxiLoadQueue.scala 131:41:@9242.4]
  wire  _T_8420; // @[AxiLoadQueue.scala 131:9:@9243.4]
  wire  storesToCheck_3_2; // @[AxiLoadQueue.scala 130:10:@9244.4]
  wire  _T_8426; // @[AxiLoadQueue.scala 130:81:@9247.4]
  wire  _T_8427; // @[AxiLoadQueue.scala 130:72:@9248.4]
  wire  _T_8429; // @[AxiLoadQueue.scala 131:33:@9249.4]
  wire  _T_8432; // @[AxiLoadQueue.scala 131:41:@9251.4]
  wire  _T_8434; // @[AxiLoadQueue.scala 131:9:@9252.4]
  wire  storesToCheck_3_3; // @[AxiLoadQueue.scala 130:10:@9253.4]
  wire  _T_8440; // @[AxiLoadQueue.scala 130:81:@9256.4]
  wire  _T_8441; // @[AxiLoadQueue.scala 130:72:@9257.4]
  wire  _T_8443; // @[AxiLoadQueue.scala 131:33:@9258.4]
  wire  _T_8446; // @[AxiLoadQueue.scala 131:41:@9260.4]
  wire  _T_8448; // @[AxiLoadQueue.scala 131:9:@9261.4]
  wire  storesToCheck_3_4; // @[AxiLoadQueue.scala 130:10:@9262.4]
  wire  _T_8454; // @[AxiLoadQueue.scala 130:81:@9265.4]
  wire  _T_8455; // @[AxiLoadQueue.scala 130:72:@9266.4]
  wire  _T_8457; // @[AxiLoadQueue.scala 131:33:@9267.4]
  wire  _T_8460; // @[AxiLoadQueue.scala 131:41:@9269.4]
  wire  _T_8462; // @[AxiLoadQueue.scala 131:9:@9270.4]
  wire  storesToCheck_3_5; // @[AxiLoadQueue.scala 130:10:@9271.4]
  wire  _T_8468; // @[AxiLoadQueue.scala 130:81:@9274.4]
  wire  _T_8469; // @[AxiLoadQueue.scala 130:72:@9275.4]
  wire  _T_8471; // @[AxiLoadQueue.scala 131:33:@9276.4]
  wire  _T_8474; // @[AxiLoadQueue.scala 131:41:@9278.4]
  wire  _T_8476; // @[AxiLoadQueue.scala 131:9:@9279.4]
  wire  storesToCheck_3_6; // @[AxiLoadQueue.scala 130:10:@9280.4]
  wire  _T_8482; // @[AxiLoadQueue.scala 130:81:@9283.4]
  wire  _T_8483; // @[AxiLoadQueue.scala 130:72:@9284.4]
  wire  _T_8485; // @[AxiLoadQueue.scala 131:33:@9285.4]
  wire  _T_8488; // @[AxiLoadQueue.scala 131:41:@9287.4]
  wire  _T_8490; // @[AxiLoadQueue.scala 131:9:@9288.4]
  wire  storesToCheck_3_7; // @[AxiLoadQueue.scala 130:10:@9289.4]
  wire  _T_8496; // @[AxiLoadQueue.scala 130:81:@9292.4]
  wire  _T_8497; // @[AxiLoadQueue.scala 130:72:@9293.4]
  wire  _T_8499; // @[AxiLoadQueue.scala 131:33:@9294.4]
  wire  _T_8502; // @[AxiLoadQueue.scala 131:41:@9296.4]
  wire  _T_8504; // @[AxiLoadQueue.scala 131:9:@9297.4]
  wire  storesToCheck_3_8; // @[AxiLoadQueue.scala 130:10:@9298.4]
  wire  _T_8510; // @[AxiLoadQueue.scala 130:81:@9301.4]
  wire  _T_8511; // @[AxiLoadQueue.scala 130:72:@9302.4]
  wire  _T_8513; // @[AxiLoadQueue.scala 131:33:@9303.4]
  wire  _T_8516; // @[AxiLoadQueue.scala 131:41:@9305.4]
  wire  _T_8518; // @[AxiLoadQueue.scala 131:9:@9306.4]
  wire  storesToCheck_3_9; // @[AxiLoadQueue.scala 130:10:@9307.4]
  wire  _T_8524; // @[AxiLoadQueue.scala 130:81:@9310.4]
  wire  _T_8525; // @[AxiLoadQueue.scala 130:72:@9311.4]
  wire  _T_8527; // @[AxiLoadQueue.scala 131:33:@9312.4]
  wire  _T_8530; // @[AxiLoadQueue.scala 131:41:@9314.4]
  wire  _T_8532; // @[AxiLoadQueue.scala 131:9:@9315.4]
  wire  storesToCheck_3_10; // @[AxiLoadQueue.scala 130:10:@9316.4]
  wire  _T_8538; // @[AxiLoadQueue.scala 130:81:@9319.4]
  wire  _T_8539; // @[AxiLoadQueue.scala 130:72:@9320.4]
  wire  _T_8541; // @[AxiLoadQueue.scala 131:33:@9321.4]
  wire  _T_8544; // @[AxiLoadQueue.scala 131:41:@9323.4]
  wire  _T_8546; // @[AxiLoadQueue.scala 131:9:@9324.4]
  wire  storesToCheck_3_11; // @[AxiLoadQueue.scala 130:10:@9325.4]
  wire  _T_8552; // @[AxiLoadQueue.scala 130:81:@9328.4]
  wire  _T_8553; // @[AxiLoadQueue.scala 130:72:@9329.4]
  wire  _T_8555; // @[AxiLoadQueue.scala 131:33:@9330.4]
  wire  _T_8558; // @[AxiLoadQueue.scala 131:41:@9332.4]
  wire  _T_8560; // @[AxiLoadQueue.scala 131:9:@9333.4]
  wire  storesToCheck_3_12; // @[AxiLoadQueue.scala 130:10:@9334.4]
  wire  _T_8566; // @[AxiLoadQueue.scala 130:81:@9337.4]
  wire  _T_8567; // @[AxiLoadQueue.scala 130:72:@9338.4]
  wire  _T_8569; // @[AxiLoadQueue.scala 131:33:@9339.4]
  wire  _T_8572; // @[AxiLoadQueue.scala 131:41:@9341.4]
  wire  _T_8574; // @[AxiLoadQueue.scala 131:9:@9342.4]
  wire  storesToCheck_3_13; // @[AxiLoadQueue.scala 130:10:@9343.4]
  wire  _T_8580; // @[AxiLoadQueue.scala 130:81:@9346.4]
  wire  _T_8581; // @[AxiLoadQueue.scala 130:72:@9347.4]
  wire  _T_8583; // @[AxiLoadQueue.scala 131:33:@9348.4]
  wire  _T_8586; // @[AxiLoadQueue.scala 131:41:@9350.4]
  wire  _T_8588; // @[AxiLoadQueue.scala 131:9:@9351.4]
  wire  storesToCheck_3_14; // @[AxiLoadQueue.scala 130:10:@9352.4]
  wire  _T_8594; // @[AxiLoadQueue.scala 130:81:@9355.4]
  wire  storesToCheck_3_15; // @[AxiLoadQueue.scala 130:10:@9361.4]
  wire  storesToCheck_4_0; // @[AxiLoadQueue.scala 130:10:@9403.4]
  wire  _T_8644; // @[AxiLoadQueue.scala 130:81:@9406.4]
  wire  _T_8645; // @[AxiLoadQueue.scala 130:72:@9407.4]
  wire  _T_8647; // @[AxiLoadQueue.scala 131:33:@9408.4]
  wire  _T_8650; // @[AxiLoadQueue.scala 131:41:@9410.4]
  wire  _T_8652; // @[AxiLoadQueue.scala 131:9:@9411.4]
  wire  storesToCheck_4_1; // @[AxiLoadQueue.scala 130:10:@9412.4]
  wire  _T_8658; // @[AxiLoadQueue.scala 130:81:@9415.4]
  wire  _T_8659; // @[AxiLoadQueue.scala 130:72:@9416.4]
  wire  _T_8661; // @[AxiLoadQueue.scala 131:33:@9417.4]
  wire  _T_8664; // @[AxiLoadQueue.scala 131:41:@9419.4]
  wire  _T_8666; // @[AxiLoadQueue.scala 131:9:@9420.4]
  wire  storesToCheck_4_2; // @[AxiLoadQueue.scala 130:10:@9421.4]
  wire  _T_8672; // @[AxiLoadQueue.scala 130:81:@9424.4]
  wire  _T_8673; // @[AxiLoadQueue.scala 130:72:@9425.4]
  wire  _T_8675; // @[AxiLoadQueue.scala 131:33:@9426.4]
  wire  _T_8678; // @[AxiLoadQueue.scala 131:41:@9428.4]
  wire  _T_8680; // @[AxiLoadQueue.scala 131:9:@9429.4]
  wire  storesToCheck_4_3; // @[AxiLoadQueue.scala 130:10:@9430.4]
  wire  _T_8686; // @[AxiLoadQueue.scala 130:81:@9433.4]
  wire  _T_8687; // @[AxiLoadQueue.scala 130:72:@9434.4]
  wire  _T_8689; // @[AxiLoadQueue.scala 131:33:@9435.4]
  wire  _T_8692; // @[AxiLoadQueue.scala 131:41:@9437.4]
  wire  _T_8694; // @[AxiLoadQueue.scala 131:9:@9438.4]
  wire  storesToCheck_4_4; // @[AxiLoadQueue.scala 130:10:@9439.4]
  wire  _T_8700; // @[AxiLoadQueue.scala 130:81:@9442.4]
  wire  _T_8701; // @[AxiLoadQueue.scala 130:72:@9443.4]
  wire  _T_8703; // @[AxiLoadQueue.scala 131:33:@9444.4]
  wire  _T_8706; // @[AxiLoadQueue.scala 131:41:@9446.4]
  wire  _T_8708; // @[AxiLoadQueue.scala 131:9:@9447.4]
  wire  storesToCheck_4_5; // @[AxiLoadQueue.scala 130:10:@9448.4]
  wire  _T_8714; // @[AxiLoadQueue.scala 130:81:@9451.4]
  wire  _T_8715; // @[AxiLoadQueue.scala 130:72:@9452.4]
  wire  _T_8717; // @[AxiLoadQueue.scala 131:33:@9453.4]
  wire  _T_8720; // @[AxiLoadQueue.scala 131:41:@9455.4]
  wire  _T_8722; // @[AxiLoadQueue.scala 131:9:@9456.4]
  wire  storesToCheck_4_6; // @[AxiLoadQueue.scala 130:10:@9457.4]
  wire  _T_8728; // @[AxiLoadQueue.scala 130:81:@9460.4]
  wire  _T_8729; // @[AxiLoadQueue.scala 130:72:@9461.4]
  wire  _T_8731; // @[AxiLoadQueue.scala 131:33:@9462.4]
  wire  _T_8734; // @[AxiLoadQueue.scala 131:41:@9464.4]
  wire  _T_8736; // @[AxiLoadQueue.scala 131:9:@9465.4]
  wire  storesToCheck_4_7; // @[AxiLoadQueue.scala 130:10:@9466.4]
  wire  _T_8742; // @[AxiLoadQueue.scala 130:81:@9469.4]
  wire  _T_8743; // @[AxiLoadQueue.scala 130:72:@9470.4]
  wire  _T_8745; // @[AxiLoadQueue.scala 131:33:@9471.4]
  wire  _T_8748; // @[AxiLoadQueue.scala 131:41:@9473.4]
  wire  _T_8750; // @[AxiLoadQueue.scala 131:9:@9474.4]
  wire  storesToCheck_4_8; // @[AxiLoadQueue.scala 130:10:@9475.4]
  wire  _T_8756; // @[AxiLoadQueue.scala 130:81:@9478.4]
  wire  _T_8757; // @[AxiLoadQueue.scala 130:72:@9479.4]
  wire  _T_8759; // @[AxiLoadQueue.scala 131:33:@9480.4]
  wire  _T_8762; // @[AxiLoadQueue.scala 131:41:@9482.4]
  wire  _T_8764; // @[AxiLoadQueue.scala 131:9:@9483.4]
  wire  storesToCheck_4_9; // @[AxiLoadQueue.scala 130:10:@9484.4]
  wire  _T_8770; // @[AxiLoadQueue.scala 130:81:@9487.4]
  wire  _T_8771; // @[AxiLoadQueue.scala 130:72:@9488.4]
  wire  _T_8773; // @[AxiLoadQueue.scala 131:33:@9489.4]
  wire  _T_8776; // @[AxiLoadQueue.scala 131:41:@9491.4]
  wire  _T_8778; // @[AxiLoadQueue.scala 131:9:@9492.4]
  wire  storesToCheck_4_10; // @[AxiLoadQueue.scala 130:10:@9493.4]
  wire  _T_8784; // @[AxiLoadQueue.scala 130:81:@9496.4]
  wire  _T_8785; // @[AxiLoadQueue.scala 130:72:@9497.4]
  wire  _T_8787; // @[AxiLoadQueue.scala 131:33:@9498.4]
  wire  _T_8790; // @[AxiLoadQueue.scala 131:41:@9500.4]
  wire  _T_8792; // @[AxiLoadQueue.scala 131:9:@9501.4]
  wire  storesToCheck_4_11; // @[AxiLoadQueue.scala 130:10:@9502.4]
  wire  _T_8798; // @[AxiLoadQueue.scala 130:81:@9505.4]
  wire  _T_8799; // @[AxiLoadQueue.scala 130:72:@9506.4]
  wire  _T_8801; // @[AxiLoadQueue.scala 131:33:@9507.4]
  wire  _T_8804; // @[AxiLoadQueue.scala 131:41:@9509.4]
  wire  _T_8806; // @[AxiLoadQueue.scala 131:9:@9510.4]
  wire  storesToCheck_4_12; // @[AxiLoadQueue.scala 130:10:@9511.4]
  wire  _T_8812; // @[AxiLoadQueue.scala 130:81:@9514.4]
  wire  _T_8813; // @[AxiLoadQueue.scala 130:72:@9515.4]
  wire  _T_8815; // @[AxiLoadQueue.scala 131:33:@9516.4]
  wire  _T_8818; // @[AxiLoadQueue.scala 131:41:@9518.4]
  wire  _T_8820; // @[AxiLoadQueue.scala 131:9:@9519.4]
  wire  storesToCheck_4_13; // @[AxiLoadQueue.scala 130:10:@9520.4]
  wire  _T_8826; // @[AxiLoadQueue.scala 130:81:@9523.4]
  wire  _T_8827; // @[AxiLoadQueue.scala 130:72:@9524.4]
  wire  _T_8829; // @[AxiLoadQueue.scala 131:33:@9525.4]
  wire  _T_8832; // @[AxiLoadQueue.scala 131:41:@9527.4]
  wire  _T_8834; // @[AxiLoadQueue.scala 131:9:@9528.4]
  wire  storesToCheck_4_14; // @[AxiLoadQueue.scala 130:10:@9529.4]
  wire  _T_8840; // @[AxiLoadQueue.scala 130:81:@9532.4]
  wire  storesToCheck_4_15; // @[AxiLoadQueue.scala 130:10:@9538.4]
  wire  storesToCheck_5_0; // @[AxiLoadQueue.scala 130:10:@9580.4]
  wire  _T_8890; // @[AxiLoadQueue.scala 130:81:@9583.4]
  wire  _T_8891; // @[AxiLoadQueue.scala 130:72:@9584.4]
  wire  _T_8893; // @[AxiLoadQueue.scala 131:33:@9585.4]
  wire  _T_8896; // @[AxiLoadQueue.scala 131:41:@9587.4]
  wire  _T_8898; // @[AxiLoadQueue.scala 131:9:@9588.4]
  wire  storesToCheck_5_1; // @[AxiLoadQueue.scala 130:10:@9589.4]
  wire  _T_8904; // @[AxiLoadQueue.scala 130:81:@9592.4]
  wire  _T_8905; // @[AxiLoadQueue.scala 130:72:@9593.4]
  wire  _T_8907; // @[AxiLoadQueue.scala 131:33:@9594.4]
  wire  _T_8910; // @[AxiLoadQueue.scala 131:41:@9596.4]
  wire  _T_8912; // @[AxiLoadQueue.scala 131:9:@9597.4]
  wire  storesToCheck_5_2; // @[AxiLoadQueue.scala 130:10:@9598.4]
  wire  _T_8918; // @[AxiLoadQueue.scala 130:81:@9601.4]
  wire  _T_8919; // @[AxiLoadQueue.scala 130:72:@9602.4]
  wire  _T_8921; // @[AxiLoadQueue.scala 131:33:@9603.4]
  wire  _T_8924; // @[AxiLoadQueue.scala 131:41:@9605.4]
  wire  _T_8926; // @[AxiLoadQueue.scala 131:9:@9606.4]
  wire  storesToCheck_5_3; // @[AxiLoadQueue.scala 130:10:@9607.4]
  wire  _T_8932; // @[AxiLoadQueue.scala 130:81:@9610.4]
  wire  _T_8933; // @[AxiLoadQueue.scala 130:72:@9611.4]
  wire  _T_8935; // @[AxiLoadQueue.scala 131:33:@9612.4]
  wire  _T_8938; // @[AxiLoadQueue.scala 131:41:@9614.4]
  wire  _T_8940; // @[AxiLoadQueue.scala 131:9:@9615.4]
  wire  storesToCheck_5_4; // @[AxiLoadQueue.scala 130:10:@9616.4]
  wire  _T_8946; // @[AxiLoadQueue.scala 130:81:@9619.4]
  wire  _T_8947; // @[AxiLoadQueue.scala 130:72:@9620.4]
  wire  _T_8949; // @[AxiLoadQueue.scala 131:33:@9621.4]
  wire  _T_8952; // @[AxiLoadQueue.scala 131:41:@9623.4]
  wire  _T_8954; // @[AxiLoadQueue.scala 131:9:@9624.4]
  wire  storesToCheck_5_5; // @[AxiLoadQueue.scala 130:10:@9625.4]
  wire  _T_8960; // @[AxiLoadQueue.scala 130:81:@9628.4]
  wire  _T_8961; // @[AxiLoadQueue.scala 130:72:@9629.4]
  wire  _T_8963; // @[AxiLoadQueue.scala 131:33:@9630.4]
  wire  _T_8966; // @[AxiLoadQueue.scala 131:41:@9632.4]
  wire  _T_8968; // @[AxiLoadQueue.scala 131:9:@9633.4]
  wire  storesToCheck_5_6; // @[AxiLoadQueue.scala 130:10:@9634.4]
  wire  _T_8974; // @[AxiLoadQueue.scala 130:81:@9637.4]
  wire  _T_8975; // @[AxiLoadQueue.scala 130:72:@9638.4]
  wire  _T_8977; // @[AxiLoadQueue.scala 131:33:@9639.4]
  wire  _T_8980; // @[AxiLoadQueue.scala 131:41:@9641.4]
  wire  _T_8982; // @[AxiLoadQueue.scala 131:9:@9642.4]
  wire  storesToCheck_5_7; // @[AxiLoadQueue.scala 130:10:@9643.4]
  wire  _T_8988; // @[AxiLoadQueue.scala 130:81:@9646.4]
  wire  _T_8989; // @[AxiLoadQueue.scala 130:72:@9647.4]
  wire  _T_8991; // @[AxiLoadQueue.scala 131:33:@9648.4]
  wire  _T_8994; // @[AxiLoadQueue.scala 131:41:@9650.4]
  wire  _T_8996; // @[AxiLoadQueue.scala 131:9:@9651.4]
  wire  storesToCheck_5_8; // @[AxiLoadQueue.scala 130:10:@9652.4]
  wire  _T_9002; // @[AxiLoadQueue.scala 130:81:@9655.4]
  wire  _T_9003; // @[AxiLoadQueue.scala 130:72:@9656.4]
  wire  _T_9005; // @[AxiLoadQueue.scala 131:33:@9657.4]
  wire  _T_9008; // @[AxiLoadQueue.scala 131:41:@9659.4]
  wire  _T_9010; // @[AxiLoadQueue.scala 131:9:@9660.4]
  wire  storesToCheck_5_9; // @[AxiLoadQueue.scala 130:10:@9661.4]
  wire  _T_9016; // @[AxiLoadQueue.scala 130:81:@9664.4]
  wire  _T_9017; // @[AxiLoadQueue.scala 130:72:@9665.4]
  wire  _T_9019; // @[AxiLoadQueue.scala 131:33:@9666.4]
  wire  _T_9022; // @[AxiLoadQueue.scala 131:41:@9668.4]
  wire  _T_9024; // @[AxiLoadQueue.scala 131:9:@9669.4]
  wire  storesToCheck_5_10; // @[AxiLoadQueue.scala 130:10:@9670.4]
  wire  _T_9030; // @[AxiLoadQueue.scala 130:81:@9673.4]
  wire  _T_9031; // @[AxiLoadQueue.scala 130:72:@9674.4]
  wire  _T_9033; // @[AxiLoadQueue.scala 131:33:@9675.4]
  wire  _T_9036; // @[AxiLoadQueue.scala 131:41:@9677.4]
  wire  _T_9038; // @[AxiLoadQueue.scala 131:9:@9678.4]
  wire  storesToCheck_5_11; // @[AxiLoadQueue.scala 130:10:@9679.4]
  wire  _T_9044; // @[AxiLoadQueue.scala 130:81:@9682.4]
  wire  _T_9045; // @[AxiLoadQueue.scala 130:72:@9683.4]
  wire  _T_9047; // @[AxiLoadQueue.scala 131:33:@9684.4]
  wire  _T_9050; // @[AxiLoadQueue.scala 131:41:@9686.4]
  wire  _T_9052; // @[AxiLoadQueue.scala 131:9:@9687.4]
  wire  storesToCheck_5_12; // @[AxiLoadQueue.scala 130:10:@9688.4]
  wire  _T_9058; // @[AxiLoadQueue.scala 130:81:@9691.4]
  wire  _T_9059; // @[AxiLoadQueue.scala 130:72:@9692.4]
  wire  _T_9061; // @[AxiLoadQueue.scala 131:33:@9693.4]
  wire  _T_9064; // @[AxiLoadQueue.scala 131:41:@9695.4]
  wire  _T_9066; // @[AxiLoadQueue.scala 131:9:@9696.4]
  wire  storesToCheck_5_13; // @[AxiLoadQueue.scala 130:10:@9697.4]
  wire  _T_9072; // @[AxiLoadQueue.scala 130:81:@9700.4]
  wire  _T_9073; // @[AxiLoadQueue.scala 130:72:@9701.4]
  wire  _T_9075; // @[AxiLoadQueue.scala 131:33:@9702.4]
  wire  _T_9078; // @[AxiLoadQueue.scala 131:41:@9704.4]
  wire  _T_9080; // @[AxiLoadQueue.scala 131:9:@9705.4]
  wire  storesToCheck_5_14; // @[AxiLoadQueue.scala 130:10:@9706.4]
  wire  _T_9086; // @[AxiLoadQueue.scala 130:81:@9709.4]
  wire  storesToCheck_5_15; // @[AxiLoadQueue.scala 130:10:@9715.4]
  wire  storesToCheck_6_0; // @[AxiLoadQueue.scala 130:10:@9757.4]
  wire  _T_9136; // @[AxiLoadQueue.scala 130:81:@9760.4]
  wire  _T_9137; // @[AxiLoadQueue.scala 130:72:@9761.4]
  wire  _T_9139; // @[AxiLoadQueue.scala 131:33:@9762.4]
  wire  _T_9142; // @[AxiLoadQueue.scala 131:41:@9764.4]
  wire  _T_9144; // @[AxiLoadQueue.scala 131:9:@9765.4]
  wire  storesToCheck_6_1; // @[AxiLoadQueue.scala 130:10:@9766.4]
  wire  _T_9150; // @[AxiLoadQueue.scala 130:81:@9769.4]
  wire  _T_9151; // @[AxiLoadQueue.scala 130:72:@9770.4]
  wire  _T_9153; // @[AxiLoadQueue.scala 131:33:@9771.4]
  wire  _T_9156; // @[AxiLoadQueue.scala 131:41:@9773.4]
  wire  _T_9158; // @[AxiLoadQueue.scala 131:9:@9774.4]
  wire  storesToCheck_6_2; // @[AxiLoadQueue.scala 130:10:@9775.4]
  wire  _T_9164; // @[AxiLoadQueue.scala 130:81:@9778.4]
  wire  _T_9165; // @[AxiLoadQueue.scala 130:72:@9779.4]
  wire  _T_9167; // @[AxiLoadQueue.scala 131:33:@9780.4]
  wire  _T_9170; // @[AxiLoadQueue.scala 131:41:@9782.4]
  wire  _T_9172; // @[AxiLoadQueue.scala 131:9:@9783.4]
  wire  storesToCheck_6_3; // @[AxiLoadQueue.scala 130:10:@9784.4]
  wire  _T_9178; // @[AxiLoadQueue.scala 130:81:@9787.4]
  wire  _T_9179; // @[AxiLoadQueue.scala 130:72:@9788.4]
  wire  _T_9181; // @[AxiLoadQueue.scala 131:33:@9789.4]
  wire  _T_9184; // @[AxiLoadQueue.scala 131:41:@9791.4]
  wire  _T_9186; // @[AxiLoadQueue.scala 131:9:@9792.4]
  wire  storesToCheck_6_4; // @[AxiLoadQueue.scala 130:10:@9793.4]
  wire  _T_9192; // @[AxiLoadQueue.scala 130:81:@9796.4]
  wire  _T_9193; // @[AxiLoadQueue.scala 130:72:@9797.4]
  wire  _T_9195; // @[AxiLoadQueue.scala 131:33:@9798.4]
  wire  _T_9198; // @[AxiLoadQueue.scala 131:41:@9800.4]
  wire  _T_9200; // @[AxiLoadQueue.scala 131:9:@9801.4]
  wire  storesToCheck_6_5; // @[AxiLoadQueue.scala 130:10:@9802.4]
  wire  _T_9206; // @[AxiLoadQueue.scala 130:81:@9805.4]
  wire  _T_9207; // @[AxiLoadQueue.scala 130:72:@9806.4]
  wire  _T_9209; // @[AxiLoadQueue.scala 131:33:@9807.4]
  wire  _T_9212; // @[AxiLoadQueue.scala 131:41:@9809.4]
  wire  _T_9214; // @[AxiLoadQueue.scala 131:9:@9810.4]
  wire  storesToCheck_6_6; // @[AxiLoadQueue.scala 130:10:@9811.4]
  wire  _T_9220; // @[AxiLoadQueue.scala 130:81:@9814.4]
  wire  _T_9221; // @[AxiLoadQueue.scala 130:72:@9815.4]
  wire  _T_9223; // @[AxiLoadQueue.scala 131:33:@9816.4]
  wire  _T_9226; // @[AxiLoadQueue.scala 131:41:@9818.4]
  wire  _T_9228; // @[AxiLoadQueue.scala 131:9:@9819.4]
  wire  storesToCheck_6_7; // @[AxiLoadQueue.scala 130:10:@9820.4]
  wire  _T_9234; // @[AxiLoadQueue.scala 130:81:@9823.4]
  wire  _T_9235; // @[AxiLoadQueue.scala 130:72:@9824.4]
  wire  _T_9237; // @[AxiLoadQueue.scala 131:33:@9825.4]
  wire  _T_9240; // @[AxiLoadQueue.scala 131:41:@9827.4]
  wire  _T_9242; // @[AxiLoadQueue.scala 131:9:@9828.4]
  wire  storesToCheck_6_8; // @[AxiLoadQueue.scala 130:10:@9829.4]
  wire  _T_9248; // @[AxiLoadQueue.scala 130:81:@9832.4]
  wire  _T_9249; // @[AxiLoadQueue.scala 130:72:@9833.4]
  wire  _T_9251; // @[AxiLoadQueue.scala 131:33:@9834.4]
  wire  _T_9254; // @[AxiLoadQueue.scala 131:41:@9836.4]
  wire  _T_9256; // @[AxiLoadQueue.scala 131:9:@9837.4]
  wire  storesToCheck_6_9; // @[AxiLoadQueue.scala 130:10:@9838.4]
  wire  _T_9262; // @[AxiLoadQueue.scala 130:81:@9841.4]
  wire  _T_9263; // @[AxiLoadQueue.scala 130:72:@9842.4]
  wire  _T_9265; // @[AxiLoadQueue.scala 131:33:@9843.4]
  wire  _T_9268; // @[AxiLoadQueue.scala 131:41:@9845.4]
  wire  _T_9270; // @[AxiLoadQueue.scala 131:9:@9846.4]
  wire  storesToCheck_6_10; // @[AxiLoadQueue.scala 130:10:@9847.4]
  wire  _T_9276; // @[AxiLoadQueue.scala 130:81:@9850.4]
  wire  _T_9277; // @[AxiLoadQueue.scala 130:72:@9851.4]
  wire  _T_9279; // @[AxiLoadQueue.scala 131:33:@9852.4]
  wire  _T_9282; // @[AxiLoadQueue.scala 131:41:@9854.4]
  wire  _T_9284; // @[AxiLoadQueue.scala 131:9:@9855.4]
  wire  storesToCheck_6_11; // @[AxiLoadQueue.scala 130:10:@9856.4]
  wire  _T_9290; // @[AxiLoadQueue.scala 130:81:@9859.4]
  wire  _T_9291; // @[AxiLoadQueue.scala 130:72:@9860.4]
  wire  _T_9293; // @[AxiLoadQueue.scala 131:33:@9861.4]
  wire  _T_9296; // @[AxiLoadQueue.scala 131:41:@9863.4]
  wire  _T_9298; // @[AxiLoadQueue.scala 131:9:@9864.4]
  wire  storesToCheck_6_12; // @[AxiLoadQueue.scala 130:10:@9865.4]
  wire  _T_9304; // @[AxiLoadQueue.scala 130:81:@9868.4]
  wire  _T_9305; // @[AxiLoadQueue.scala 130:72:@9869.4]
  wire  _T_9307; // @[AxiLoadQueue.scala 131:33:@9870.4]
  wire  _T_9310; // @[AxiLoadQueue.scala 131:41:@9872.4]
  wire  _T_9312; // @[AxiLoadQueue.scala 131:9:@9873.4]
  wire  storesToCheck_6_13; // @[AxiLoadQueue.scala 130:10:@9874.4]
  wire  _T_9318; // @[AxiLoadQueue.scala 130:81:@9877.4]
  wire  _T_9319; // @[AxiLoadQueue.scala 130:72:@9878.4]
  wire  _T_9321; // @[AxiLoadQueue.scala 131:33:@9879.4]
  wire  _T_9324; // @[AxiLoadQueue.scala 131:41:@9881.4]
  wire  _T_9326; // @[AxiLoadQueue.scala 131:9:@9882.4]
  wire  storesToCheck_6_14; // @[AxiLoadQueue.scala 130:10:@9883.4]
  wire  _T_9332; // @[AxiLoadQueue.scala 130:81:@9886.4]
  wire  storesToCheck_6_15; // @[AxiLoadQueue.scala 130:10:@9892.4]
  wire  storesToCheck_7_0; // @[AxiLoadQueue.scala 130:10:@9934.4]
  wire  _T_9382; // @[AxiLoadQueue.scala 130:81:@9937.4]
  wire  _T_9383; // @[AxiLoadQueue.scala 130:72:@9938.4]
  wire  _T_9385; // @[AxiLoadQueue.scala 131:33:@9939.4]
  wire  _T_9388; // @[AxiLoadQueue.scala 131:41:@9941.4]
  wire  _T_9390; // @[AxiLoadQueue.scala 131:9:@9942.4]
  wire  storesToCheck_7_1; // @[AxiLoadQueue.scala 130:10:@9943.4]
  wire  _T_9396; // @[AxiLoadQueue.scala 130:81:@9946.4]
  wire  _T_9397; // @[AxiLoadQueue.scala 130:72:@9947.4]
  wire  _T_9399; // @[AxiLoadQueue.scala 131:33:@9948.4]
  wire  _T_9402; // @[AxiLoadQueue.scala 131:41:@9950.4]
  wire  _T_9404; // @[AxiLoadQueue.scala 131:9:@9951.4]
  wire  storesToCheck_7_2; // @[AxiLoadQueue.scala 130:10:@9952.4]
  wire  _T_9410; // @[AxiLoadQueue.scala 130:81:@9955.4]
  wire  _T_9411; // @[AxiLoadQueue.scala 130:72:@9956.4]
  wire  _T_9413; // @[AxiLoadQueue.scala 131:33:@9957.4]
  wire  _T_9416; // @[AxiLoadQueue.scala 131:41:@9959.4]
  wire  _T_9418; // @[AxiLoadQueue.scala 131:9:@9960.4]
  wire  storesToCheck_7_3; // @[AxiLoadQueue.scala 130:10:@9961.4]
  wire  _T_9424; // @[AxiLoadQueue.scala 130:81:@9964.4]
  wire  _T_9425; // @[AxiLoadQueue.scala 130:72:@9965.4]
  wire  _T_9427; // @[AxiLoadQueue.scala 131:33:@9966.4]
  wire  _T_9430; // @[AxiLoadQueue.scala 131:41:@9968.4]
  wire  _T_9432; // @[AxiLoadQueue.scala 131:9:@9969.4]
  wire  storesToCheck_7_4; // @[AxiLoadQueue.scala 130:10:@9970.4]
  wire  _T_9438; // @[AxiLoadQueue.scala 130:81:@9973.4]
  wire  _T_9439; // @[AxiLoadQueue.scala 130:72:@9974.4]
  wire  _T_9441; // @[AxiLoadQueue.scala 131:33:@9975.4]
  wire  _T_9444; // @[AxiLoadQueue.scala 131:41:@9977.4]
  wire  _T_9446; // @[AxiLoadQueue.scala 131:9:@9978.4]
  wire  storesToCheck_7_5; // @[AxiLoadQueue.scala 130:10:@9979.4]
  wire  _T_9452; // @[AxiLoadQueue.scala 130:81:@9982.4]
  wire  _T_9453; // @[AxiLoadQueue.scala 130:72:@9983.4]
  wire  _T_9455; // @[AxiLoadQueue.scala 131:33:@9984.4]
  wire  _T_9458; // @[AxiLoadQueue.scala 131:41:@9986.4]
  wire  _T_9460; // @[AxiLoadQueue.scala 131:9:@9987.4]
  wire  storesToCheck_7_6; // @[AxiLoadQueue.scala 130:10:@9988.4]
  wire  _T_9466; // @[AxiLoadQueue.scala 130:81:@9991.4]
  wire  _T_9467; // @[AxiLoadQueue.scala 130:72:@9992.4]
  wire  _T_9469; // @[AxiLoadQueue.scala 131:33:@9993.4]
  wire  _T_9472; // @[AxiLoadQueue.scala 131:41:@9995.4]
  wire  _T_9474; // @[AxiLoadQueue.scala 131:9:@9996.4]
  wire  storesToCheck_7_7; // @[AxiLoadQueue.scala 130:10:@9997.4]
  wire  _T_9480; // @[AxiLoadQueue.scala 130:81:@10000.4]
  wire  _T_9481; // @[AxiLoadQueue.scala 130:72:@10001.4]
  wire  _T_9483; // @[AxiLoadQueue.scala 131:33:@10002.4]
  wire  _T_9486; // @[AxiLoadQueue.scala 131:41:@10004.4]
  wire  _T_9488; // @[AxiLoadQueue.scala 131:9:@10005.4]
  wire  storesToCheck_7_8; // @[AxiLoadQueue.scala 130:10:@10006.4]
  wire  _T_9494; // @[AxiLoadQueue.scala 130:81:@10009.4]
  wire  _T_9495; // @[AxiLoadQueue.scala 130:72:@10010.4]
  wire  _T_9497; // @[AxiLoadQueue.scala 131:33:@10011.4]
  wire  _T_9500; // @[AxiLoadQueue.scala 131:41:@10013.4]
  wire  _T_9502; // @[AxiLoadQueue.scala 131:9:@10014.4]
  wire  storesToCheck_7_9; // @[AxiLoadQueue.scala 130:10:@10015.4]
  wire  _T_9508; // @[AxiLoadQueue.scala 130:81:@10018.4]
  wire  _T_9509; // @[AxiLoadQueue.scala 130:72:@10019.4]
  wire  _T_9511; // @[AxiLoadQueue.scala 131:33:@10020.4]
  wire  _T_9514; // @[AxiLoadQueue.scala 131:41:@10022.4]
  wire  _T_9516; // @[AxiLoadQueue.scala 131:9:@10023.4]
  wire  storesToCheck_7_10; // @[AxiLoadQueue.scala 130:10:@10024.4]
  wire  _T_9522; // @[AxiLoadQueue.scala 130:81:@10027.4]
  wire  _T_9523; // @[AxiLoadQueue.scala 130:72:@10028.4]
  wire  _T_9525; // @[AxiLoadQueue.scala 131:33:@10029.4]
  wire  _T_9528; // @[AxiLoadQueue.scala 131:41:@10031.4]
  wire  _T_9530; // @[AxiLoadQueue.scala 131:9:@10032.4]
  wire  storesToCheck_7_11; // @[AxiLoadQueue.scala 130:10:@10033.4]
  wire  _T_9536; // @[AxiLoadQueue.scala 130:81:@10036.4]
  wire  _T_9537; // @[AxiLoadQueue.scala 130:72:@10037.4]
  wire  _T_9539; // @[AxiLoadQueue.scala 131:33:@10038.4]
  wire  _T_9542; // @[AxiLoadQueue.scala 131:41:@10040.4]
  wire  _T_9544; // @[AxiLoadQueue.scala 131:9:@10041.4]
  wire  storesToCheck_7_12; // @[AxiLoadQueue.scala 130:10:@10042.4]
  wire  _T_9550; // @[AxiLoadQueue.scala 130:81:@10045.4]
  wire  _T_9551; // @[AxiLoadQueue.scala 130:72:@10046.4]
  wire  _T_9553; // @[AxiLoadQueue.scala 131:33:@10047.4]
  wire  _T_9556; // @[AxiLoadQueue.scala 131:41:@10049.4]
  wire  _T_9558; // @[AxiLoadQueue.scala 131:9:@10050.4]
  wire  storesToCheck_7_13; // @[AxiLoadQueue.scala 130:10:@10051.4]
  wire  _T_9564; // @[AxiLoadQueue.scala 130:81:@10054.4]
  wire  _T_9565; // @[AxiLoadQueue.scala 130:72:@10055.4]
  wire  _T_9567; // @[AxiLoadQueue.scala 131:33:@10056.4]
  wire  _T_9570; // @[AxiLoadQueue.scala 131:41:@10058.4]
  wire  _T_9572; // @[AxiLoadQueue.scala 131:9:@10059.4]
  wire  storesToCheck_7_14; // @[AxiLoadQueue.scala 130:10:@10060.4]
  wire  _T_9578; // @[AxiLoadQueue.scala 130:81:@10063.4]
  wire  storesToCheck_7_15; // @[AxiLoadQueue.scala 130:10:@10069.4]
  wire  storesToCheck_8_0; // @[AxiLoadQueue.scala 130:10:@10111.4]
  wire  _T_9628; // @[AxiLoadQueue.scala 130:81:@10114.4]
  wire  _T_9629; // @[AxiLoadQueue.scala 130:72:@10115.4]
  wire  _T_9631; // @[AxiLoadQueue.scala 131:33:@10116.4]
  wire  _T_9634; // @[AxiLoadQueue.scala 131:41:@10118.4]
  wire  _T_9636; // @[AxiLoadQueue.scala 131:9:@10119.4]
  wire  storesToCheck_8_1; // @[AxiLoadQueue.scala 130:10:@10120.4]
  wire  _T_9642; // @[AxiLoadQueue.scala 130:81:@10123.4]
  wire  _T_9643; // @[AxiLoadQueue.scala 130:72:@10124.4]
  wire  _T_9645; // @[AxiLoadQueue.scala 131:33:@10125.4]
  wire  _T_9648; // @[AxiLoadQueue.scala 131:41:@10127.4]
  wire  _T_9650; // @[AxiLoadQueue.scala 131:9:@10128.4]
  wire  storesToCheck_8_2; // @[AxiLoadQueue.scala 130:10:@10129.4]
  wire  _T_9656; // @[AxiLoadQueue.scala 130:81:@10132.4]
  wire  _T_9657; // @[AxiLoadQueue.scala 130:72:@10133.4]
  wire  _T_9659; // @[AxiLoadQueue.scala 131:33:@10134.4]
  wire  _T_9662; // @[AxiLoadQueue.scala 131:41:@10136.4]
  wire  _T_9664; // @[AxiLoadQueue.scala 131:9:@10137.4]
  wire  storesToCheck_8_3; // @[AxiLoadQueue.scala 130:10:@10138.4]
  wire  _T_9670; // @[AxiLoadQueue.scala 130:81:@10141.4]
  wire  _T_9671; // @[AxiLoadQueue.scala 130:72:@10142.4]
  wire  _T_9673; // @[AxiLoadQueue.scala 131:33:@10143.4]
  wire  _T_9676; // @[AxiLoadQueue.scala 131:41:@10145.4]
  wire  _T_9678; // @[AxiLoadQueue.scala 131:9:@10146.4]
  wire  storesToCheck_8_4; // @[AxiLoadQueue.scala 130:10:@10147.4]
  wire  _T_9684; // @[AxiLoadQueue.scala 130:81:@10150.4]
  wire  _T_9685; // @[AxiLoadQueue.scala 130:72:@10151.4]
  wire  _T_9687; // @[AxiLoadQueue.scala 131:33:@10152.4]
  wire  _T_9690; // @[AxiLoadQueue.scala 131:41:@10154.4]
  wire  _T_9692; // @[AxiLoadQueue.scala 131:9:@10155.4]
  wire  storesToCheck_8_5; // @[AxiLoadQueue.scala 130:10:@10156.4]
  wire  _T_9698; // @[AxiLoadQueue.scala 130:81:@10159.4]
  wire  _T_9699; // @[AxiLoadQueue.scala 130:72:@10160.4]
  wire  _T_9701; // @[AxiLoadQueue.scala 131:33:@10161.4]
  wire  _T_9704; // @[AxiLoadQueue.scala 131:41:@10163.4]
  wire  _T_9706; // @[AxiLoadQueue.scala 131:9:@10164.4]
  wire  storesToCheck_8_6; // @[AxiLoadQueue.scala 130:10:@10165.4]
  wire  _T_9712; // @[AxiLoadQueue.scala 130:81:@10168.4]
  wire  _T_9713; // @[AxiLoadQueue.scala 130:72:@10169.4]
  wire  _T_9715; // @[AxiLoadQueue.scala 131:33:@10170.4]
  wire  _T_9718; // @[AxiLoadQueue.scala 131:41:@10172.4]
  wire  _T_9720; // @[AxiLoadQueue.scala 131:9:@10173.4]
  wire  storesToCheck_8_7; // @[AxiLoadQueue.scala 130:10:@10174.4]
  wire  _T_9726; // @[AxiLoadQueue.scala 130:81:@10177.4]
  wire  _T_9727; // @[AxiLoadQueue.scala 130:72:@10178.4]
  wire  _T_9729; // @[AxiLoadQueue.scala 131:33:@10179.4]
  wire  _T_9732; // @[AxiLoadQueue.scala 131:41:@10181.4]
  wire  _T_9734; // @[AxiLoadQueue.scala 131:9:@10182.4]
  wire  storesToCheck_8_8; // @[AxiLoadQueue.scala 130:10:@10183.4]
  wire  _T_9740; // @[AxiLoadQueue.scala 130:81:@10186.4]
  wire  _T_9741; // @[AxiLoadQueue.scala 130:72:@10187.4]
  wire  _T_9743; // @[AxiLoadQueue.scala 131:33:@10188.4]
  wire  _T_9746; // @[AxiLoadQueue.scala 131:41:@10190.4]
  wire  _T_9748; // @[AxiLoadQueue.scala 131:9:@10191.4]
  wire  storesToCheck_8_9; // @[AxiLoadQueue.scala 130:10:@10192.4]
  wire  _T_9754; // @[AxiLoadQueue.scala 130:81:@10195.4]
  wire  _T_9755; // @[AxiLoadQueue.scala 130:72:@10196.4]
  wire  _T_9757; // @[AxiLoadQueue.scala 131:33:@10197.4]
  wire  _T_9760; // @[AxiLoadQueue.scala 131:41:@10199.4]
  wire  _T_9762; // @[AxiLoadQueue.scala 131:9:@10200.4]
  wire  storesToCheck_8_10; // @[AxiLoadQueue.scala 130:10:@10201.4]
  wire  _T_9768; // @[AxiLoadQueue.scala 130:81:@10204.4]
  wire  _T_9769; // @[AxiLoadQueue.scala 130:72:@10205.4]
  wire  _T_9771; // @[AxiLoadQueue.scala 131:33:@10206.4]
  wire  _T_9774; // @[AxiLoadQueue.scala 131:41:@10208.4]
  wire  _T_9776; // @[AxiLoadQueue.scala 131:9:@10209.4]
  wire  storesToCheck_8_11; // @[AxiLoadQueue.scala 130:10:@10210.4]
  wire  _T_9782; // @[AxiLoadQueue.scala 130:81:@10213.4]
  wire  _T_9783; // @[AxiLoadQueue.scala 130:72:@10214.4]
  wire  _T_9785; // @[AxiLoadQueue.scala 131:33:@10215.4]
  wire  _T_9788; // @[AxiLoadQueue.scala 131:41:@10217.4]
  wire  _T_9790; // @[AxiLoadQueue.scala 131:9:@10218.4]
  wire  storesToCheck_8_12; // @[AxiLoadQueue.scala 130:10:@10219.4]
  wire  _T_9796; // @[AxiLoadQueue.scala 130:81:@10222.4]
  wire  _T_9797; // @[AxiLoadQueue.scala 130:72:@10223.4]
  wire  _T_9799; // @[AxiLoadQueue.scala 131:33:@10224.4]
  wire  _T_9802; // @[AxiLoadQueue.scala 131:41:@10226.4]
  wire  _T_9804; // @[AxiLoadQueue.scala 131:9:@10227.4]
  wire  storesToCheck_8_13; // @[AxiLoadQueue.scala 130:10:@10228.4]
  wire  _T_9810; // @[AxiLoadQueue.scala 130:81:@10231.4]
  wire  _T_9811; // @[AxiLoadQueue.scala 130:72:@10232.4]
  wire  _T_9813; // @[AxiLoadQueue.scala 131:33:@10233.4]
  wire  _T_9816; // @[AxiLoadQueue.scala 131:41:@10235.4]
  wire  _T_9818; // @[AxiLoadQueue.scala 131:9:@10236.4]
  wire  storesToCheck_8_14; // @[AxiLoadQueue.scala 130:10:@10237.4]
  wire  _T_9824; // @[AxiLoadQueue.scala 130:81:@10240.4]
  wire  storesToCheck_8_15; // @[AxiLoadQueue.scala 130:10:@10246.4]
  wire  storesToCheck_9_0; // @[AxiLoadQueue.scala 130:10:@10288.4]
  wire  _T_9874; // @[AxiLoadQueue.scala 130:81:@10291.4]
  wire  _T_9875; // @[AxiLoadQueue.scala 130:72:@10292.4]
  wire  _T_9877; // @[AxiLoadQueue.scala 131:33:@10293.4]
  wire  _T_9880; // @[AxiLoadQueue.scala 131:41:@10295.4]
  wire  _T_9882; // @[AxiLoadQueue.scala 131:9:@10296.4]
  wire  storesToCheck_9_1; // @[AxiLoadQueue.scala 130:10:@10297.4]
  wire  _T_9888; // @[AxiLoadQueue.scala 130:81:@10300.4]
  wire  _T_9889; // @[AxiLoadQueue.scala 130:72:@10301.4]
  wire  _T_9891; // @[AxiLoadQueue.scala 131:33:@10302.4]
  wire  _T_9894; // @[AxiLoadQueue.scala 131:41:@10304.4]
  wire  _T_9896; // @[AxiLoadQueue.scala 131:9:@10305.4]
  wire  storesToCheck_9_2; // @[AxiLoadQueue.scala 130:10:@10306.4]
  wire  _T_9902; // @[AxiLoadQueue.scala 130:81:@10309.4]
  wire  _T_9903; // @[AxiLoadQueue.scala 130:72:@10310.4]
  wire  _T_9905; // @[AxiLoadQueue.scala 131:33:@10311.4]
  wire  _T_9908; // @[AxiLoadQueue.scala 131:41:@10313.4]
  wire  _T_9910; // @[AxiLoadQueue.scala 131:9:@10314.4]
  wire  storesToCheck_9_3; // @[AxiLoadQueue.scala 130:10:@10315.4]
  wire  _T_9916; // @[AxiLoadQueue.scala 130:81:@10318.4]
  wire  _T_9917; // @[AxiLoadQueue.scala 130:72:@10319.4]
  wire  _T_9919; // @[AxiLoadQueue.scala 131:33:@10320.4]
  wire  _T_9922; // @[AxiLoadQueue.scala 131:41:@10322.4]
  wire  _T_9924; // @[AxiLoadQueue.scala 131:9:@10323.4]
  wire  storesToCheck_9_4; // @[AxiLoadQueue.scala 130:10:@10324.4]
  wire  _T_9930; // @[AxiLoadQueue.scala 130:81:@10327.4]
  wire  _T_9931; // @[AxiLoadQueue.scala 130:72:@10328.4]
  wire  _T_9933; // @[AxiLoadQueue.scala 131:33:@10329.4]
  wire  _T_9936; // @[AxiLoadQueue.scala 131:41:@10331.4]
  wire  _T_9938; // @[AxiLoadQueue.scala 131:9:@10332.4]
  wire  storesToCheck_9_5; // @[AxiLoadQueue.scala 130:10:@10333.4]
  wire  _T_9944; // @[AxiLoadQueue.scala 130:81:@10336.4]
  wire  _T_9945; // @[AxiLoadQueue.scala 130:72:@10337.4]
  wire  _T_9947; // @[AxiLoadQueue.scala 131:33:@10338.4]
  wire  _T_9950; // @[AxiLoadQueue.scala 131:41:@10340.4]
  wire  _T_9952; // @[AxiLoadQueue.scala 131:9:@10341.4]
  wire  storesToCheck_9_6; // @[AxiLoadQueue.scala 130:10:@10342.4]
  wire  _T_9958; // @[AxiLoadQueue.scala 130:81:@10345.4]
  wire  _T_9959; // @[AxiLoadQueue.scala 130:72:@10346.4]
  wire  _T_9961; // @[AxiLoadQueue.scala 131:33:@10347.4]
  wire  _T_9964; // @[AxiLoadQueue.scala 131:41:@10349.4]
  wire  _T_9966; // @[AxiLoadQueue.scala 131:9:@10350.4]
  wire  storesToCheck_9_7; // @[AxiLoadQueue.scala 130:10:@10351.4]
  wire  _T_9972; // @[AxiLoadQueue.scala 130:81:@10354.4]
  wire  _T_9973; // @[AxiLoadQueue.scala 130:72:@10355.4]
  wire  _T_9975; // @[AxiLoadQueue.scala 131:33:@10356.4]
  wire  _T_9978; // @[AxiLoadQueue.scala 131:41:@10358.4]
  wire  _T_9980; // @[AxiLoadQueue.scala 131:9:@10359.4]
  wire  storesToCheck_9_8; // @[AxiLoadQueue.scala 130:10:@10360.4]
  wire  _T_9986; // @[AxiLoadQueue.scala 130:81:@10363.4]
  wire  _T_9987; // @[AxiLoadQueue.scala 130:72:@10364.4]
  wire  _T_9989; // @[AxiLoadQueue.scala 131:33:@10365.4]
  wire  _T_9992; // @[AxiLoadQueue.scala 131:41:@10367.4]
  wire  _T_9994; // @[AxiLoadQueue.scala 131:9:@10368.4]
  wire  storesToCheck_9_9; // @[AxiLoadQueue.scala 130:10:@10369.4]
  wire  _T_10000; // @[AxiLoadQueue.scala 130:81:@10372.4]
  wire  _T_10001; // @[AxiLoadQueue.scala 130:72:@10373.4]
  wire  _T_10003; // @[AxiLoadQueue.scala 131:33:@10374.4]
  wire  _T_10006; // @[AxiLoadQueue.scala 131:41:@10376.4]
  wire  _T_10008; // @[AxiLoadQueue.scala 131:9:@10377.4]
  wire  storesToCheck_9_10; // @[AxiLoadQueue.scala 130:10:@10378.4]
  wire  _T_10014; // @[AxiLoadQueue.scala 130:81:@10381.4]
  wire  _T_10015; // @[AxiLoadQueue.scala 130:72:@10382.4]
  wire  _T_10017; // @[AxiLoadQueue.scala 131:33:@10383.4]
  wire  _T_10020; // @[AxiLoadQueue.scala 131:41:@10385.4]
  wire  _T_10022; // @[AxiLoadQueue.scala 131:9:@10386.4]
  wire  storesToCheck_9_11; // @[AxiLoadQueue.scala 130:10:@10387.4]
  wire  _T_10028; // @[AxiLoadQueue.scala 130:81:@10390.4]
  wire  _T_10029; // @[AxiLoadQueue.scala 130:72:@10391.4]
  wire  _T_10031; // @[AxiLoadQueue.scala 131:33:@10392.4]
  wire  _T_10034; // @[AxiLoadQueue.scala 131:41:@10394.4]
  wire  _T_10036; // @[AxiLoadQueue.scala 131:9:@10395.4]
  wire  storesToCheck_9_12; // @[AxiLoadQueue.scala 130:10:@10396.4]
  wire  _T_10042; // @[AxiLoadQueue.scala 130:81:@10399.4]
  wire  _T_10043; // @[AxiLoadQueue.scala 130:72:@10400.4]
  wire  _T_10045; // @[AxiLoadQueue.scala 131:33:@10401.4]
  wire  _T_10048; // @[AxiLoadQueue.scala 131:41:@10403.4]
  wire  _T_10050; // @[AxiLoadQueue.scala 131:9:@10404.4]
  wire  storesToCheck_9_13; // @[AxiLoadQueue.scala 130:10:@10405.4]
  wire  _T_10056; // @[AxiLoadQueue.scala 130:81:@10408.4]
  wire  _T_10057; // @[AxiLoadQueue.scala 130:72:@10409.4]
  wire  _T_10059; // @[AxiLoadQueue.scala 131:33:@10410.4]
  wire  _T_10062; // @[AxiLoadQueue.scala 131:41:@10412.4]
  wire  _T_10064; // @[AxiLoadQueue.scala 131:9:@10413.4]
  wire  storesToCheck_9_14; // @[AxiLoadQueue.scala 130:10:@10414.4]
  wire  _T_10070; // @[AxiLoadQueue.scala 130:81:@10417.4]
  wire  storesToCheck_9_15; // @[AxiLoadQueue.scala 130:10:@10423.4]
  wire  storesToCheck_10_0; // @[AxiLoadQueue.scala 130:10:@10465.4]
  wire  _T_10120; // @[AxiLoadQueue.scala 130:81:@10468.4]
  wire  _T_10121; // @[AxiLoadQueue.scala 130:72:@10469.4]
  wire  _T_10123; // @[AxiLoadQueue.scala 131:33:@10470.4]
  wire  _T_10126; // @[AxiLoadQueue.scala 131:41:@10472.4]
  wire  _T_10128; // @[AxiLoadQueue.scala 131:9:@10473.4]
  wire  storesToCheck_10_1; // @[AxiLoadQueue.scala 130:10:@10474.4]
  wire  _T_10134; // @[AxiLoadQueue.scala 130:81:@10477.4]
  wire  _T_10135; // @[AxiLoadQueue.scala 130:72:@10478.4]
  wire  _T_10137; // @[AxiLoadQueue.scala 131:33:@10479.4]
  wire  _T_10140; // @[AxiLoadQueue.scala 131:41:@10481.4]
  wire  _T_10142; // @[AxiLoadQueue.scala 131:9:@10482.4]
  wire  storesToCheck_10_2; // @[AxiLoadQueue.scala 130:10:@10483.4]
  wire  _T_10148; // @[AxiLoadQueue.scala 130:81:@10486.4]
  wire  _T_10149; // @[AxiLoadQueue.scala 130:72:@10487.4]
  wire  _T_10151; // @[AxiLoadQueue.scala 131:33:@10488.4]
  wire  _T_10154; // @[AxiLoadQueue.scala 131:41:@10490.4]
  wire  _T_10156; // @[AxiLoadQueue.scala 131:9:@10491.4]
  wire  storesToCheck_10_3; // @[AxiLoadQueue.scala 130:10:@10492.4]
  wire  _T_10162; // @[AxiLoadQueue.scala 130:81:@10495.4]
  wire  _T_10163; // @[AxiLoadQueue.scala 130:72:@10496.4]
  wire  _T_10165; // @[AxiLoadQueue.scala 131:33:@10497.4]
  wire  _T_10168; // @[AxiLoadQueue.scala 131:41:@10499.4]
  wire  _T_10170; // @[AxiLoadQueue.scala 131:9:@10500.4]
  wire  storesToCheck_10_4; // @[AxiLoadQueue.scala 130:10:@10501.4]
  wire  _T_10176; // @[AxiLoadQueue.scala 130:81:@10504.4]
  wire  _T_10177; // @[AxiLoadQueue.scala 130:72:@10505.4]
  wire  _T_10179; // @[AxiLoadQueue.scala 131:33:@10506.4]
  wire  _T_10182; // @[AxiLoadQueue.scala 131:41:@10508.4]
  wire  _T_10184; // @[AxiLoadQueue.scala 131:9:@10509.4]
  wire  storesToCheck_10_5; // @[AxiLoadQueue.scala 130:10:@10510.4]
  wire  _T_10190; // @[AxiLoadQueue.scala 130:81:@10513.4]
  wire  _T_10191; // @[AxiLoadQueue.scala 130:72:@10514.4]
  wire  _T_10193; // @[AxiLoadQueue.scala 131:33:@10515.4]
  wire  _T_10196; // @[AxiLoadQueue.scala 131:41:@10517.4]
  wire  _T_10198; // @[AxiLoadQueue.scala 131:9:@10518.4]
  wire  storesToCheck_10_6; // @[AxiLoadQueue.scala 130:10:@10519.4]
  wire  _T_10204; // @[AxiLoadQueue.scala 130:81:@10522.4]
  wire  _T_10205; // @[AxiLoadQueue.scala 130:72:@10523.4]
  wire  _T_10207; // @[AxiLoadQueue.scala 131:33:@10524.4]
  wire  _T_10210; // @[AxiLoadQueue.scala 131:41:@10526.4]
  wire  _T_10212; // @[AxiLoadQueue.scala 131:9:@10527.4]
  wire  storesToCheck_10_7; // @[AxiLoadQueue.scala 130:10:@10528.4]
  wire  _T_10218; // @[AxiLoadQueue.scala 130:81:@10531.4]
  wire  _T_10219; // @[AxiLoadQueue.scala 130:72:@10532.4]
  wire  _T_10221; // @[AxiLoadQueue.scala 131:33:@10533.4]
  wire  _T_10224; // @[AxiLoadQueue.scala 131:41:@10535.4]
  wire  _T_10226; // @[AxiLoadQueue.scala 131:9:@10536.4]
  wire  storesToCheck_10_8; // @[AxiLoadQueue.scala 130:10:@10537.4]
  wire  _T_10232; // @[AxiLoadQueue.scala 130:81:@10540.4]
  wire  _T_10233; // @[AxiLoadQueue.scala 130:72:@10541.4]
  wire  _T_10235; // @[AxiLoadQueue.scala 131:33:@10542.4]
  wire  _T_10238; // @[AxiLoadQueue.scala 131:41:@10544.4]
  wire  _T_10240; // @[AxiLoadQueue.scala 131:9:@10545.4]
  wire  storesToCheck_10_9; // @[AxiLoadQueue.scala 130:10:@10546.4]
  wire  _T_10246; // @[AxiLoadQueue.scala 130:81:@10549.4]
  wire  _T_10247; // @[AxiLoadQueue.scala 130:72:@10550.4]
  wire  _T_10249; // @[AxiLoadQueue.scala 131:33:@10551.4]
  wire  _T_10252; // @[AxiLoadQueue.scala 131:41:@10553.4]
  wire  _T_10254; // @[AxiLoadQueue.scala 131:9:@10554.4]
  wire  storesToCheck_10_10; // @[AxiLoadQueue.scala 130:10:@10555.4]
  wire  _T_10260; // @[AxiLoadQueue.scala 130:81:@10558.4]
  wire  _T_10261; // @[AxiLoadQueue.scala 130:72:@10559.4]
  wire  _T_10263; // @[AxiLoadQueue.scala 131:33:@10560.4]
  wire  _T_10266; // @[AxiLoadQueue.scala 131:41:@10562.4]
  wire  _T_10268; // @[AxiLoadQueue.scala 131:9:@10563.4]
  wire  storesToCheck_10_11; // @[AxiLoadQueue.scala 130:10:@10564.4]
  wire  _T_10274; // @[AxiLoadQueue.scala 130:81:@10567.4]
  wire  _T_10275; // @[AxiLoadQueue.scala 130:72:@10568.4]
  wire  _T_10277; // @[AxiLoadQueue.scala 131:33:@10569.4]
  wire  _T_10280; // @[AxiLoadQueue.scala 131:41:@10571.4]
  wire  _T_10282; // @[AxiLoadQueue.scala 131:9:@10572.4]
  wire  storesToCheck_10_12; // @[AxiLoadQueue.scala 130:10:@10573.4]
  wire  _T_10288; // @[AxiLoadQueue.scala 130:81:@10576.4]
  wire  _T_10289; // @[AxiLoadQueue.scala 130:72:@10577.4]
  wire  _T_10291; // @[AxiLoadQueue.scala 131:33:@10578.4]
  wire  _T_10294; // @[AxiLoadQueue.scala 131:41:@10580.4]
  wire  _T_10296; // @[AxiLoadQueue.scala 131:9:@10581.4]
  wire  storesToCheck_10_13; // @[AxiLoadQueue.scala 130:10:@10582.4]
  wire  _T_10302; // @[AxiLoadQueue.scala 130:81:@10585.4]
  wire  _T_10303; // @[AxiLoadQueue.scala 130:72:@10586.4]
  wire  _T_10305; // @[AxiLoadQueue.scala 131:33:@10587.4]
  wire  _T_10308; // @[AxiLoadQueue.scala 131:41:@10589.4]
  wire  _T_10310; // @[AxiLoadQueue.scala 131:9:@10590.4]
  wire  storesToCheck_10_14; // @[AxiLoadQueue.scala 130:10:@10591.4]
  wire  _T_10316; // @[AxiLoadQueue.scala 130:81:@10594.4]
  wire  storesToCheck_10_15; // @[AxiLoadQueue.scala 130:10:@10600.4]
  wire  storesToCheck_11_0; // @[AxiLoadQueue.scala 130:10:@10642.4]
  wire  _T_10366; // @[AxiLoadQueue.scala 130:81:@10645.4]
  wire  _T_10367; // @[AxiLoadQueue.scala 130:72:@10646.4]
  wire  _T_10369; // @[AxiLoadQueue.scala 131:33:@10647.4]
  wire  _T_10372; // @[AxiLoadQueue.scala 131:41:@10649.4]
  wire  _T_10374; // @[AxiLoadQueue.scala 131:9:@10650.4]
  wire  storesToCheck_11_1; // @[AxiLoadQueue.scala 130:10:@10651.4]
  wire  _T_10380; // @[AxiLoadQueue.scala 130:81:@10654.4]
  wire  _T_10381; // @[AxiLoadQueue.scala 130:72:@10655.4]
  wire  _T_10383; // @[AxiLoadQueue.scala 131:33:@10656.4]
  wire  _T_10386; // @[AxiLoadQueue.scala 131:41:@10658.4]
  wire  _T_10388; // @[AxiLoadQueue.scala 131:9:@10659.4]
  wire  storesToCheck_11_2; // @[AxiLoadQueue.scala 130:10:@10660.4]
  wire  _T_10394; // @[AxiLoadQueue.scala 130:81:@10663.4]
  wire  _T_10395; // @[AxiLoadQueue.scala 130:72:@10664.4]
  wire  _T_10397; // @[AxiLoadQueue.scala 131:33:@10665.4]
  wire  _T_10400; // @[AxiLoadQueue.scala 131:41:@10667.4]
  wire  _T_10402; // @[AxiLoadQueue.scala 131:9:@10668.4]
  wire  storesToCheck_11_3; // @[AxiLoadQueue.scala 130:10:@10669.4]
  wire  _T_10408; // @[AxiLoadQueue.scala 130:81:@10672.4]
  wire  _T_10409; // @[AxiLoadQueue.scala 130:72:@10673.4]
  wire  _T_10411; // @[AxiLoadQueue.scala 131:33:@10674.4]
  wire  _T_10414; // @[AxiLoadQueue.scala 131:41:@10676.4]
  wire  _T_10416; // @[AxiLoadQueue.scala 131:9:@10677.4]
  wire  storesToCheck_11_4; // @[AxiLoadQueue.scala 130:10:@10678.4]
  wire  _T_10422; // @[AxiLoadQueue.scala 130:81:@10681.4]
  wire  _T_10423; // @[AxiLoadQueue.scala 130:72:@10682.4]
  wire  _T_10425; // @[AxiLoadQueue.scala 131:33:@10683.4]
  wire  _T_10428; // @[AxiLoadQueue.scala 131:41:@10685.4]
  wire  _T_10430; // @[AxiLoadQueue.scala 131:9:@10686.4]
  wire  storesToCheck_11_5; // @[AxiLoadQueue.scala 130:10:@10687.4]
  wire  _T_10436; // @[AxiLoadQueue.scala 130:81:@10690.4]
  wire  _T_10437; // @[AxiLoadQueue.scala 130:72:@10691.4]
  wire  _T_10439; // @[AxiLoadQueue.scala 131:33:@10692.4]
  wire  _T_10442; // @[AxiLoadQueue.scala 131:41:@10694.4]
  wire  _T_10444; // @[AxiLoadQueue.scala 131:9:@10695.4]
  wire  storesToCheck_11_6; // @[AxiLoadQueue.scala 130:10:@10696.4]
  wire  _T_10450; // @[AxiLoadQueue.scala 130:81:@10699.4]
  wire  _T_10451; // @[AxiLoadQueue.scala 130:72:@10700.4]
  wire  _T_10453; // @[AxiLoadQueue.scala 131:33:@10701.4]
  wire  _T_10456; // @[AxiLoadQueue.scala 131:41:@10703.4]
  wire  _T_10458; // @[AxiLoadQueue.scala 131:9:@10704.4]
  wire  storesToCheck_11_7; // @[AxiLoadQueue.scala 130:10:@10705.4]
  wire  _T_10464; // @[AxiLoadQueue.scala 130:81:@10708.4]
  wire  _T_10465; // @[AxiLoadQueue.scala 130:72:@10709.4]
  wire  _T_10467; // @[AxiLoadQueue.scala 131:33:@10710.4]
  wire  _T_10470; // @[AxiLoadQueue.scala 131:41:@10712.4]
  wire  _T_10472; // @[AxiLoadQueue.scala 131:9:@10713.4]
  wire  storesToCheck_11_8; // @[AxiLoadQueue.scala 130:10:@10714.4]
  wire  _T_10478; // @[AxiLoadQueue.scala 130:81:@10717.4]
  wire  _T_10479; // @[AxiLoadQueue.scala 130:72:@10718.4]
  wire  _T_10481; // @[AxiLoadQueue.scala 131:33:@10719.4]
  wire  _T_10484; // @[AxiLoadQueue.scala 131:41:@10721.4]
  wire  _T_10486; // @[AxiLoadQueue.scala 131:9:@10722.4]
  wire  storesToCheck_11_9; // @[AxiLoadQueue.scala 130:10:@10723.4]
  wire  _T_10492; // @[AxiLoadQueue.scala 130:81:@10726.4]
  wire  _T_10493; // @[AxiLoadQueue.scala 130:72:@10727.4]
  wire  _T_10495; // @[AxiLoadQueue.scala 131:33:@10728.4]
  wire  _T_10498; // @[AxiLoadQueue.scala 131:41:@10730.4]
  wire  _T_10500; // @[AxiLoadQueue.scala 131:9:@10731.4]
  wire  storesToCheck_11_10; // @[AxiLoadQueue.scala 130:10:@10732.4]
  wire  _T_10506; // @[AxiLoadQueue.scala 130:81:@10735.4]
  wire  _T_10507; // @[AxiLoadQueue.scala 130:72:@10736.4]
  wire  _T_10509; // @[AxiLoadQueue.scala 131:33:@10737.4]
  wire  _T_10512; // @[AxiLoadQueue.scala 131:41:@10739.4]
  wire  _T_10514; // @[AxiLoadQueue.scala 131:9:@10740.4]
  wire  storesToCheck_11_11; // @[AxiLoadQueue.scala 130:10:@10741.4]
  wire  _T_10520; // @[AxiLoadQueue.scala 130:81:@10744.4]
  wire  _T_10521; // @[AxiLoadQueue.scala 130:72:@10745.4]
  wire  _T_10523; // @[AxiLoadQueue.scala 131:33:@10746.4]
  wire  _T_10526; // @[AxiLoadQueue.scala 131:41:@10748.4]
  wire  _T_10528; // @[AxiLoadQueue.scala 131:9:@10749.4]
  wire  storesToCheck_11_12; // @[AxiLoadQueue.scala 130:10:@10750.4]
  wire  _T_10534; // @[AxiLoadQueue.scala 130:81:@10753.4]
  wire  _T_10535; // @[AxiLoadQueue.scala 130:72:@10754.4]
  wire  _T_10537; // @[AxiLoadQueue.scala 131:33:@10755.4]
  wire  _T_10540; // @[AxiLoadQueue.scala 131:41:@10757.4]
  wire  _T_10542; // @[AxiLoadQueue.scala 131:9:@10758.4]
  wire  storesToCheck_11_13; // @[AxiLoadQueue.scala 130:10:@10759.4]
  wire  _T_10548; // @[AxiLoadQueue.scala 130:81:@10762.4]
  wire  _T_10549; // @[AxiLoadQueue.scala 130:72:@10763.4]
  wire  _T_10551; // @[AxiLoadQueue.scala 131:33:@10764.4]
  wire  _T_10554; // @[AxiLoadQueue.scala 131:41:@10766.4]
  wire  _T_10556; // @[AxiLoadQueue.scala 131:9:@10767.4]
  wire  storesToCheck_11_14; // @[AxiLoadQueue.scala 130:10:@10768.4]
  wire  _T_10562; // @[AxiLoadQueue.scala 130:81:@10771.4]
  wire  storesToCheck_11_15; // @[AxiLoadQueue.scala 130:10:@10777.4]
  wire  storesToCheck_12_0; // @[AxiLoadQueue.scala 130:10:@10819.4]
  wire  _T_10612; // @[AxiLoadQueue.scala 130:81:@10822.4]
  wire  _T_10613; // @[AxiLoadQueue.scala 130:72:@10823.4]
  wire  _T_10615; // @[AxiLoadQueue.scala 131:33:@10824.4]
  wire  _T_10618; // @[AxiLoadQueue.scala 131:41:@10826.4]
  wire  _T_10620; // @[AxiLoadQueue.scala 131:9:@10827.4]
  wire  storesToCheck_12_1; // @[AxiLoadQueue.scala 130:10:@10828.4]
  wire  _T_10626; // @[AxiLoadQueue.scala 130:81:@10831.4]
  wire  _T_10627; // @[AxiLoadQueue.scala 130:72:@10832.4]
  wire  _T_10629; // @[AxiLoadQueue.scala 131:33:@10833.4]
  wire  _T_10632; // @[AxiLoadQueue.scala 131:41:@10835.4]
  wire  _T_10634; // @[AxiLoadQueue.scala 131:9:@10836.4]
  wire  storesToCheck_12_2; // @[AxiLoadQueue.scala 130:10:@10837.4]
  wire  _T_10640; // @[AxiLoadQueue.scala 130:81:@10840.4]
  wire  _T_10641; // @[AxiLoadQueue.scala 130:72:@10841.4]
  wire  _T_10643; // @[AxiLoadQueue.scala 131:33:@10842.4]
  wire  _T_10646; // @[AxiLoadQueue.scala 131:41:@10844.4]
  wire  _T_10648; // @[AxiLoadQueue.scala 131:9:@10845.4]
  wire  storesToCheck_12_3; // @[AxiLoadQueue.scala 130:10:@10846.4]
  wire  _T_10654; // @[AxiLoadQueue.scala 130:81:@10849.4]
  wire  _T_10655; // @[AxiLoadQueue.scala 130:72:@10850.4]
  wire  _T_10657; // @[AxiLoadQueue.scala 131:33:@10851.4]
  wire  _T_10660; // @[AxiLoadQueue.scala 131:41:@10853.4]
  wire  _T_10662; // @[AxiLoadQueue.scala 131:9:@10854.4]
  wire  storesToCheck_12_4; // @[AxiLoadQueue.scala 130:10:@10855.4]
  wire  _T_10668; // @[AxiLoadQueue.scala 130:81:@10858.4]
  wire  _T_10669; // @[AxiLoadQueue.scala 130:72:@10859.4]
  wire  _T_10671; // @[AxiLoadQueue.scala 131:33:@10860.4]
  wire  _T_10674; // @[AxiLoadQueue.scala 131:41:@10862.4]
  wire  _T_10676; // @[AxiLoadQueue.scala 131:9:@10863.4]
  wire  storesToCheck_12_5; // @[AxiLoadQueue.scala 130:10:@10864.4]
  wire  _T_10682; // @[AxiLoadQueue.scala 130:81:@10867.4]
  wire  _T_10683; // @[AxiLoadQueue.scala 130:72:@10868.4]
  wire  _T_10685; // @[AxiLoadQueue.scala 131:33:@10869.4]
  wire  _T_10688; // @[AxiLoadQueue.scala 131:41:@10871.4]
  wire  _T_10690; // @[AxiLoadQueue.scala 131:9:@10872.4]
  wire  storesToCheck_12_6; // @[AxiLoadQueue.scala 130:10:@10873.4]
  wire  _T_10696; // @[AxiLoadQueue.scala 130:81:@10876.4]
  wire  _T_10697; // @[AxiLoadQueue.scala 130:72:@10877.4]
  wire  _T_10699; // @[AxiLoadQueue.scala 131:33:@10878.4]
  wire  _T_10702; // @[AxiLoadQueue.scala 131:41:@10880.4]
  wire  _T_10704; // @[AxiLoadQueue.scala 131:9:@10881.4]
  wire  storesToCheck_12_7; // @[AxiLoadQueue.scala 130:10:@10882.4]
  wire  _T_10710; // @[AxiLoadQueue.scala 130:81:@10885.4]
  wire  _T_10711; // @[AxiLoadQueue.scala 130:72:@10886.4]
  wire  _T_10713; // @[AxiLoadQueue.scala 131:33:@10887.4]
  wire  _T_10716; // @[AxiLoadQueue.scala 131:41:@10889.4]
  wire  _T_10718; // @[AxiLoadQueue.scala 131:9:@10890.4]
  wire  storesToCheck_12_8; // @[AxiLoadQueue.scala 130:10:@10891.4]
  wire  _T_10724; // @[AxiLoadQueue.scala 130:81:@10894.4]
  wire  _T_10725; // @[AxiLoadQueue.scala 130:72:@10895.4]
  wire  _T_10727; // @[AxiLoadQueue.scala 131:33:@10896.4]
  wire  _T_10730; // @[AxiLoadQueue.scala 131:41:@10898.4]
  wire  _T_10732; // @[AxiLoadQueue.scala 131:9:@10899.4]
  wire  storesToCheck_12_9; // @[AxiLoadQueue.scala 130:10:@10900.4]
  wire  _T_10738; // @[AxiLoadQueue.scala 130:81:@10903.4]
  wire  _T_10739; // @[AxiLoadQueue.scala 130:72:@10904.4]
  wire  _T_10741; // @[AxiLoadQueue.scala 131:33:@10905.4]
  wire  _T_10744; // @[AxiLoadQueue.scala 131:41:@10907.4]
  wire  _T_10746; // @[AxiLoadQueue.scala 131:9:@10908.4]
  wire  storesToCheck_12_10; // @[AxiLoadQueue.scala 130:10:@10909.4]
  wire  _T_10752; // @[AxiLoadQueue.scala 130:81:@10912.4]
  wire  _T_10753; // @[AxiLoadQueue.scala 130:72:@10913.4]
  wire  _T_10755; // @[AxiLoadQueue.scala 131:33:@10914.4]
  wire  _T_10758; // @[AxiLoadQueue.scala 131:41:@10916.4]
  wire  _T_10760; // @[AxiLoadQueue.scala 131:9:@10917.4]
  wire  storesToCheck_12_11; // @[AxiLoadQueue.scala 130:10:@10918.4]
  wire  _T_10766; // @[AxiLoadQueue.scala 130:81:@10921.4]
  wire  _T_10767; // @[AxiLoadQueue.scala 130:72:@10922.4]
  wire  _T_10769; // @[AxiLoadQueue.scala 131:33:@10923.4]
  wire  _T_10772; // @[AxiLoadQueue.scala 131:41:@10925.4]
  wire  _T_10774; // @[AxiLoadQueue.scala 131:9:@10926.4]
  wire  storesToCheck_12_12; // @[AxiLoadQueue.scala 130:10:@10927.4]
  wire  _T_10780; // @[AxiLoadQueue.scala 130:81:@10930.4]
  wire  _T_10781; // @[AxiLoadQueue.scala 130:72:@10931.4]
  wire  _T_10783; // @[AxiLoadQueue.scala 131:33:@10932.4]
  wire  _T_10786; // @[AxiLoadQueue.scala 131:41:@10934.4]
  wire  _T_10788; // @[AxiLoadQueue.scala 131:9:@10935.4]
  wire  storesToCheck_12_13; // @[AxiLoadQueue.scala 130:10:@10936.4]
  wire  _T_10794; // @[AxiLoadQueue.scala 130:81:@10939.4]
  wire  _T_10795; // @[AxiLoadQueue.scala 130:72:@10940.4]
  wire  _T_10797; // @[AxiLoadQueue.scala 131:33:@10941.4]
  wire  _T_10800; // @[AxiLoadQueue.scala 131:41:@10943.4]
  wire  _T_10802; // @[AxiLoadQueue.scala 131:9:@10944.4]
  wire  storesToCheck_12_14; // @[AxiLoadQueue.scala 130:10:@10945.4]
  wire  _T_10808; // @[AxiLoadQueue.scala 130:81:@10948.4]
  wire  storesToCheck_12_15; // @[AxiLoadQueue.scala 130:10:@10954.4]
  wire  storesToCheck_13_0; // @[AxiLoadQueue.scala 130:10:@10996.4]
  wire  _T_10858; // @[AxiLoadQueue.scala 130:81:@10999.4]
  wire  _T_10859; // @[AxiLoadQueue.scala 130:72:@11000.4]
  wire  _T_10861; // @[AxiLoadQueue.scala 131:33:@11001.4]
  wire  _T_10864; // @[AxiLoadQueue.scala 131:41:@11003.4]
  wire  _T_10866; // @[AxiLoadQueue.scala 131:9:@11004.4]
  wire  storesToCheck_13_1; // @[AxiLoadQueue.scala 130:10:@11005.4]
  wire  _T_10872; // @[AxiLoadQueue.scala 130:81:@11008.4]
  wire  _T_10873; // @[AxiLoadQueue.scala 130:72:@11009.4]
  wire  _T_10875; // @[AxiLoadQueue.scala 131:33:@11010.4]
  wire  _T_10878; // @[AxiLoadQueue.scala 131:41:@11012.4]
  wire  _T_10880; // @[AxiLoadQueue.scala 131:9:@11013.4]
  wire  storesToCheck_13_2; // @[AxiLoadQueue.scala 130:10:@11014.4]
  wire  _T_10886; // @[AxiLoadQueue.scala 130:81:@11017.4]
  wire  _T_10887; // @[AxiLoadQueue.scala 130:72:@11018.4]
  wire  _T_10889; // @[AxiLoadQueue.scala 131:33:@11019.4]
  wire  _T_10892; // @[AxiLoadQueue.scala 131:41:@11021.4]
  wire  _T_10894; // @[AxiLoadQueue.scala 131:9:@11022.4]
  wire  storesToCheck_13_3; // @[AxiLoadQueue.scala 130:10:@11023.4]
  wire  _T_10900; // @[AxiLoadQueue.scala 130:81:@11026.4]
  wire  _T_10901; // @[AxiLoadQueue.scala 130:72:@11027.4]
  wire  _T_10903; // @[AxiLoadQueue.scala 131:33:@11028.4]
  wire  _T_10906; // @[AxiLoadQueue.scala 131:41:@11030.4]
  wire  _T_10908; // @[AxiLoadQueue.scala 131:9:@11031.4]
  wire  storesToCheck_13_4; // @[AxiLoadQueue.scala 130:10:@11032.4]
  wire  _T_10914; // @[AxiLoadQueue.scala 130:81:@11035.4]
  wire  _T_10915; // @[AxiLoadQueue.scala 130:72:@11036.4]
  wire  _T_10917; // @[AxiLoadQueue.scala 131:33:@11037.4]
  wire  _T_10920; // @[AxiLoadQueue.scala 131:41:@11039.4]
  wire  _T_10922; // @[AxiLoadQueue.scala 131:9:@11040.4]
  wire  storesToCheck_13_5; // @[AxiLoadQueue.scala 130:10:@11041.4]
  wire  _T_10928; // @[AxiLoadQueue.scala 130:81:@11044.4]
  wire  _T_10929; // @[AxiLoadQueue.scala 130:72:@11045.4]
  wire  _T_10931; // @[AxiLoadQueue.scala 131:33:@11046.4]
  wire  _T_10934; // @[AxiLoadQueue.scala 131:41:@11048.4]
  wire  _T_10936; // @[AxiLoadQueue.scala 131:9:@11049.4]
  wire  storesToCheck_13_6; // @[AxiLoadQueue.scala 130:10:@11050.4]
  wire  _T_10942; // @[AxiLoadQueue.scala 130:81:@11053.4]
  wire  _T_10943; // @[AxiLoadQueue.scala 130:72:@11054.4]
  wire  _T_10945; // @[AxiLoadQueue.scala 131:33:@11055.4]
  wire  _T_10948; // @[AxiLoadQueue.scala 131:41:@11057.4]
  wire  _T_10950; // @[AxiLoadQueue.scala 131:9:@11058.4]
  wire  storesToCheck_13_7; // @[AxiLoadQueue.scala 130:10:@11059.4]
  wire  _T_10956; // @[AxiLoadQueue.scala 130:81:@11062.4]
  wire  _T_10957; // @[AxiLoadQueue.scala 130:72:@11063.4]
  wire  _T_10959; // @[AxiLoadQueue.scala 131:33:@11064.4]
  wire  _T_10962; // @[AxiLoadQueue.scala 131:41:@11066.4]
  wire  _T_10964; // @[AxiLoadQueue.scala 131:9:@11067.4]
  wire  storesToCheck_13_8; // @[AxiLoadQueue.scala 130:10:@11068.4]
  wire  _T_10970; // @[AxiLoadQueue.scala 130:81:@11071.4]
  wire  _T_10971; // @[AxiLoadQueue.scala 130:72:@11072.4]
  wire  _T_10973; // @[AxiLoadQueue.scala 131:33:@11073.4]
  wire  _T_10976; // @[AxiLoadQueue.scala 131:41:@11075.4]
  wire  _T_10978; // @[AxiLoadQueue.scala 131:9:@11076.4]
  wire  storesToCheck_13_9; // @[AxiLoadQueue.scala 130:10:@11077.4]
  wire  _T_10984; // @[AxiLoadQueue.scala 130:81:@11080.4]
  wire  _T_10985; // @[AxiLoadQueue.scala 130:72:@11081.4]
  wire  _T_10987; // @[AxiLoadQueue.scala 131:33:@11082.4]
  wire  _T_10990; // @[AxiLoadQueue.scala 131:41:@11084.4]
  wire  _T_10992; // @[AxiLoadQueue.scala 131:9:@11085.4]
  wire  storesToCheck_13_10; // @[AxiLoadQueue.scala 130:10:@11086.4]
  wire  _T_10998; // @[AxiLoadQueue.scala 130:81:@11089.4]
  wire  _T_10999; // @[AxiLoadQueue.scala 130:72:@11090.4]
  wire  _T_11001; // @[AxiLoadQueue.scala 131:33:@11091.4]
  wire  _T_11004; // @[AxiLoadQueue.scala 131:41:@11093.4]
  wire  _T_11006; // @[AxiLoadQueue.scala 131:9:@11094.4]
  wire  storesToCheck_13_11; // @[AxiLoadQueue.scala 130:10:@11095.4]
  wire  _T_11012; // @[AxiLoadQueue.scala 130:81:@11098.4]
  wire  _T_11013; // @[AxiLoadQueue.scala 130:72:@11099.4]
  wire  _T_11015; // @[AxiLoadQueue.scala 131:33:@11100.4]
  wire  _T_11018; // @[AxiLoadQueue.scala 131:41:@11102.4]
  wire  _T_11020; // @[AxiLoadQueue.scala 131:9:@11103.4]
  wire  storesToCheck_13_12; // @[AxiLoadQueue.scala 130:10:@11104.4]
  wire  _T_11026; // @[AxiLoadQueue.scala 130:81:@11107.4]
  wire  _T_11027; // @[AxiLoadQueue.scala 130:72:@11108.4]
  wire  _T_11029; // @[AxiLoadQueue.scala 131:33:@11109.4]
  wire  _T_11032; // @[AxiLoadQueue.scala 131:41:@11111.4]
  wire  _T_11034; // @[AxiLoadQueue.scala 131:9:@11112.4]
  wire  storesToCheck_13_13; // @[AxiLoadQueue.scala 130:10:@11113.4]
  wire  _T_11040; // @[AxiLoadQueue.scala 130:81:@11116.4]
  wire  _T_11041; // @[AxiLoadQueue.scala 130:72:@11117.4]
  wire  _T_11043; // @[AxiLoadQueue.scala 131:33:@11118.4]
  wire  _T_11046; // @[AxiLoadQueue.scala 131:41:@11120.4]
  wire  _T_11048; // @[AxiLoadQueue.scala 131:9:@11121.4]
  wire  storesToCheck_13_14; // @[AxiLoadQueue.scala 130:10:@11122.4]
  wire  _T_11054; // @[AxiLoadQueue.scala 130:81:@11125.4]
  wire  storesToCheck_13_15; // @[AxiLoadQueue.scala 130:10:@11131.4]
  wire  storesToCheck_14_0; // @[AxiLoadQueue.scala 130:10:@11173.4]
  wire  _T_11104; // @[AxiLoadQueue.scala 130:81:@11176.4]
  wire  _T_11105; // @[AxiLoadQueue.scala 130:72:@11177.4]
  wire  _T_11107; // @[AxiLoadQueue.scala 131:33:@11178.4]
  wire  _T_11110; // @[AxiLoadQueue.scala 131:41:@11180.4]
  wire  _T_11112; // @[AxiLoadQueue.scala 131:9:@11181.4]
  wire  storesToCheck_14_1; // @[AxiLoadQueue.scala 130:10:@11182.4]
  wire  _T_11118; // @[AxiLoadQueue.scala 130:81:@11185.4]
  wire  _T_11119; // @[AxiLoadQueue.scala 130:72:@11186.4]
  wire  _T_11121; // @[AxiLoadQueue.scala 131:33:@11187.4]
  wire  _T_11124; // @[AxiLoadQueue.scala 131:41:@11189.4]
  wire  _T_11126; // @[AxiLoadQueue.scala 131:9:@11190.4]
  wire  storesToCheck_14_2; // @[AxiLoadQueue.scala 130:10:@11191.4]
  wire  _T_11132; // @[AxiLoadQueue.scala 130:81:@11194.4]
  wire  _T_11133; // @[AxiLoadQueue.scala 130:72:@11195.4]
  wire  _T_11135; // @[AxiLoadQueue.scala 131:33:@11196.4]
  wire  _T_11138; // @[AxiLoadQueue.scala 131:41:@11198.4]
  wire  _T_11140; // @[AxiLoadQueue.scala 131:9:@11199.4]
  wire  storesToCheck_14_3; // @[AxiLoadQueue.scala 130:10:@11200.4]
  wire  _T_11146; // @[AxiLoadQueue.scala 130:81:@11203.4]
  wire  _T_11147; // @[AxiLoadQueue.scala 130:72:@11204.4]
  wire  _T_11149; // @[AxiLoadQueue.scala 131:33:@11205.4]
  wire  _T_11152; // @[AxiLoadQueue.scala 131:41:@11207.4]
  wire  _T_11154; // @[AxiLoadQueue.scala 131:9:@11208.4]
  wire  storesToCheck_14_4; // @[AxiLoadQueue.scala 130:10:@11209.4]
  wire  _T_11160; // @[AxiLoadQueue.scala 130:81:@11212.4]
  wire  _T_11161; // @[AxiLoadQueue.scala 130:72:@11213.4]
  wire  _T_11163; // @[AxiLoadQueue.scala 131:33:@11214.4]
  wire  _T_11166; // @[AxiLoadQueue.scala 131:41:@11216.4]
  wire  _T_11168; // @[AxiLoadQueue.scala 131:9:@11217.4]
  wire  storesToCheck_14_5; // @[AxiLoadQueue.scala 130:10:@11218.4]
  wire  _T_11174; // @[AxiLoadQueue.scala 130:81:@11221.4]
  wire  _T_11175; // @[AxiLoadQueue.scala 130:72:@11222.4]
  wire  _T_11177; // @[AxiLoadQueue.scala 131:33:@11223.4]
  wire  _T_11180; // @[AxiLoadQueue.scala 131:41:@11225.4]
  wire  _T_11182; // @[AxiLoadQueue.scala 131:9:@11226.4]
  wire  storesToCheck_14_6; // @[AxiLoadQueue.scala 130:10:@11227.4]
  wire  _T_11188; // @[AxiLoadQueue.scala 130:81:@11230.4]
  wire  _T_11189; // @[AxiLoadQueue.scala 130:72:@11231.4]
  wire  _T_11191; // @[AxiLoadQueue.scala 131:33:@11232.4]
  wire  _T_11194; // @[AxiLoadQueue.scala 131:41:@11234.4]
  wire  _T_11196; // @[AxiLoadQueue.scala 131:9:@11235.4]
  wire  storesToCheck_14_7; // @[AxiLoadQueue.scala 130:10:@11236.4]
  wire  _T_11202; // @[AxiLoadQueue.scala 130:81:@11239.4]
  wire  _T_11203; // @[AxiLoadQueue.scala 130:72:@11240.4]
  wire  _T_11205; // @[AxiLoadQueue.scala 131:33:@11241.4]
  wire  _T_11208; // @[AxiLoadQueue.scala 131:41:@11243.4]
  wire  _T_11210; // @[AxiLoadQueue.scala 131:9:@11244.4]
  wire  storesToCheck_14_8; // @[AxiLoadQueue.scala 130:10:@11245.4]
  wire  _T_11216; // @[AxiLoadQueue.scala 130:81:@11248.4]
  wire  _T_11217; // @[AxiLoadQueue.scala 130:72:@11249.4]
  wire  _T_11219; // @[AxiLoadQueue.scala 131:33:@11250.4]
  wire  _T_11222; // @[AxiLoadQueue.scala 131:41:@11252.4]
  wire  _T_11224; // @[AxiLoadQueue.scala 131:9:@11253.4]
  wire  storesToCheck_14_9; // @[AxiLoadQueue.scala 130:10:@11254.4]
  wire  _T_11230; // @[AxiLoadQueue.scala 130:81:@11257.4]
  wire  _T_11231; // @[AxiLoadQueue.scala 130:72:@11258.4]
  wire  _T_11233; // @[AxiLoadQueue.scala 131:33:@11259.4]
  wire  _T_11236; // @[AxiLoadQueue.scala 131:41:@11261.4]
  wire  _T_11238; // @[AxiLoadQueue.scala 131:9:@11262.4]
  wire  storesToCheck_14_10; // @[AxiLoadQueue.scala 130:10:@11263.4]
  wire  _T_11244; // @[AxiLoadQueue.scala 130:81:@11266.4]
  wire  _T_11245; // @[AxiLoadQueue.scala 130:72:@11267.4]
  wire  _T_11247; // @[AxiLoadQueue.scala 131:33:@11268.4]
  wire  _T_11250; // @[AxiLoadQueue.scala 131:41:@11270.4]
  wire  _T_11252; // @[AxiLoadQueue.scala 131:9:@11271.4]
  wire  storesToCheck_14_11; // @[AxiLoadQueue.scala 130:10:@11272.4]
  wire  _T_11258; // @[AxiLoadQueue.scala 130:81:@11275.4]
  wire  _T_11259; // @[AxiLoadQueue.scala 130:72:@11276.4]
  wire  _T_11261; // @[AxiLoadQueue.scala 131:33:@11277.4]
  wire  _T_11264; // @[AxiLoadQueue.scala 131:41:@11279.4]
  wire  _T_11266; // @[AxiLoadQueue.scala 131:9:@11280.4]
  wire  storesToCheck_14_12; // @[AxiLoadQueue.scala 130:10:@11281.4]
  wire  _T_11272; // @[AxiLoadQueue.scala 130:81:@11284.4]
  wire  _T_11273; // @[AxiLoadQueue.scala 130:72:@11285.4]
  wire  _T_11275; // @[AxiLoadQueue.scala 131:33:@11286.4]
  wire  _T_11278; // @[AxiLoadQueue.scala 131:41:@11288.4]
  wire  _T_11280; // @[AxiLoadQueue.scala 131:9:@11289.4]
  wire  storesToCheck_14_13; // @[AxiLoadQueue.scala 130:10:@11290.4]
  wire  _T_11286; // @[AxiLoadQueue.scala 130:81:@11293.4]
  wire  _T_11287; // @[AxiLoadQueue.scala 130:72:@11294.4]
  wire  _T_11289; // @[AxiLoadQueue.scala 131:33:@11295.4]
  wire  _T_11292; // @[AxiLoadQueue.scala 131:41:@11297.4]
  wire  _T_11294; // @[AxiLoadQueue.scala 131:9:@11298.4]
  wire  storesToCheck_14_14; // @[AxiLoadQueue.scala 130:10:@11299.4]
  wire  _T_11300; // @[AxiLoadQueue.scala 130:81:@11302.4]
  wire  storesToCheck_14_15; // @[AxiLoadQueue.scala 130:10:@11308.4]
  wire  storesToCheck_15_0; // @[AxiLoadQueue.scala 130:10:@11350.4]
  wire  _T_11350; // @[AxiLoadQueue.scala 130:81:@11353.4]
  wire  _T_11351; // @[AxiLoadQueue.scala 130:72:@11354.4]
  wire  _T_11353; // @[AxiLoadQueue.scala 131:33:@11355.4]
  wire  _T_11356; // @[AxiLoadQueue.scala 131:41:@11357.4]
  wire  _T_11358; // @[AxiLoadQueue.scala 131:9:@11358.4]
  wire  storesToCheck_15_1; // @[AxiLoadQueue.scala 130:10:@11359.4]
  wire  _T_11364; // @[AxiLoadQueue.scala 130:81:@11362.4]
  wire  _T_11365; // @[AxiLoadQueue.scala 130:72:@11363.4]
  wire  _T_11367; // @[AxiLoadQueue.scala 131:33:@11364.4]
  wire  _T_11370; // @[AxiLoadQueue.scala 131:41:@11366.4]
  wire  _T_11372; // @[AxiLoadQueue.scala 131:9:@11367.4]
  wire  storesToCheck_15_2; // @[AxiLoadQueue.scala 130:10:@11368.4]
  wire  _T_11378; // @[AxiLoadQueue.scala 130:81:@11371.4]
  wire  _T_11379; // @[AxiLoadQueue.scala 130:72:@11372.4]
  wire  _T_11381; // @[AxiLoadQueue.scala 131:33:@11373.4]
  wire  _T_11384; // @[AxiLoadQueue.scala 131:41:@11375.4]
  wire  _T_11386; // @[AxiLoadQueue.scala 131:9:@11376.4]
  wire  storesToCheck_15_3; // @[AxiLoadQueue.scala 130:10:@11377.4]
  wire  _T_11392; // @[AxiLoadQueue.scala 130:81:@11380.4]
  wire  _T_11393; // @[AxiLoadQueue.scala 130:72:@11381.4]
  wire  _T_11395; // @[AxiLoadQueue.scala 131:33:@11382.4]
  wire  _T_11398; // @[AxiLoadQueue.scala 131:41:@11384.4]
  wire  _T_11400; // @[AxiLoadQueue.scala 131:9:@11385.4]
  wire  storesToCheck_15_4; // @[AxiLoadQueue.scala 130:10:@11386.4]
  wire  _T_11406; // @[AxiLoadQueue.scala 130:81:@11389.4]
  wire  _T_11407; // @[AxiLoadQueue.scala 130:72:@11390.4]
  wire  _T_11409; // @[AxiLoadQueue.scala 131:33:@11391.4]
  wire  _T_11412; // @[AxiLoadQueue.scala 131:41:@11393.4]
  wire  _T_11414; // @[AxiLoadQueue.scala 131:9:@11394.4]
  wire  storesToCheck_15_5; // @[AxiLoadQueue.scala 130:10:@11395.4]
  wire  _T_11420; // @[AxiLoadQueue.scala 130:81:@11398.4]
  wire  _T_11421; // @[AxiLoadQueue.scala 130:72:@11399.4]
  wire  _T_11423; // @[AxiLoadQueue.scala 131:33:@11400.4]
  wire  _T_11426; // @[AxiLoadQueue.scala 131:41:@11402.4]
  wire  _T_11428; // @[AxiLoadQueue.scala 131:9:@11403.4]
  wire  storesToCheck_15_6; // @[AxiLoadQueue.scala 130:10:@11404.4]
  wire  _T_11434; // @[AxiLoadQueue.scala 130:81:@11407.4]
  wire  _T_11435; // @[AxiLoadQueue.scala 130:72:@11408.4]
  wire  _T_11437; // @[AxiLoadQueue.scala 131:33:@11409.4]
  wire  _T_11440; // @[AxiLoadQueue.scala 131:41:@11411.4]
  wire  _T_11442; // @[AxiLoadQueue.scala 131:9:@11412.4]
  wire  storesToCheck_15_7; // @[AxiLoadQueue.scala 130:10:@11413.4]
  wire  _T_11448; // @[AxiLoadQueue.scala 130:81:@11416.4]
  wire  _T_11449; // @[AxiLoadQueue.scala 130:72:@11417.4]
  wire  _T_11451; // @[AxiLoadQueue.scala 131:33:@11418.4]
  wire  _T_11454; // @[AxiLoadQueue.scala 131:41:@11420.4]
  wire  _T_11456; // @[AxiLoadQueue.scala 131:9:@11421.4]
  wire  storesToCheck_15_8; // @[AxiLoadQueue.scala 130:10:@11422.4]
  wire  _T_11462; // @[AxiLoadQueue.scala 130:81:@11425.4]
  wire  _T_11463; // @[AxiLoadQueue.scala 130:72:@11426.4]
  wire  _T_11465; // @[AxiLoadQueue.scala 131:33:@11427.4]
  wire  _T_11468; // @[AxiLoadQueue.scala 131:41:@11429.4]
  wire  _T_11470; // @[AxiLoadQueue.scala 131:9:@11430.4]
  wire  storesToCheck_15_9; // @[AxiLoadQueue.scala 130:10:@11431.4]
  wire  _T_11476; // @[AxiLoadQueue.scala 130:81:@11434.4]
  wire  _T_11477; // @[AxiLoadQueue.scala 130:72:@11435.4]
  wire  _T_11479; // @[AxiLoadQueue.scala 131:33:@11436.4]
  wire  _T_11482; // @[AxiLoadQueue.scala 131:41:@11438.4]
  wire  _T_11484; // @[AxiLoadQueue.scala 131:9:@11439.4]
  wire  storesToCheck_15_10; // @[AxiLoadQueue.scala 130:10:@11440.4]
  wire  _T_11490; // @[AxiLoadQueue.scala 130:81:@11443.4]
  wire  _T_11491; // @[AxiLoadQueue.scala 130:72:@11444.4]
  wire  _T_11493; // @[AxiLoadQueue.scala 131:33:@11445.4]
  wire  _T_11496; // @[AxiLoadQueue.scala 131:41:@11447.4]
  wire  _T_11498; // @[AxiLoadQueue.scala 131:9:@11448.4]
  wire  storesToCheck_15_11; // @[AxiLoadQueue.scala 130:10:@11449.4]
  wire  _T_11504; // @[AxiLoadQueue.scala 130:81:@11452.4]
  wire  _T_11505; // @[AxiLoadQueue.scala 130:72:@11453.4]
  wire  _T_11507; // @[AxiLoadQueue.scala 131:33:@11454.4]
  wire  _T_11510; // @[AxiLoadQueue.scala 131:41:@11456.4]
  wire  _T_11512; // @[AxiLoadQueue.scala 131:9:@11457.4]
  wire  storesToCheck_15_12; // @[AxiLoadQueue.scala 130:10:@11458.4]
  wire  _T_11518; // @[AxiLoadQueue.scala 130:81:@11461.4]
  wire  _T_11519; // @[AxiLoadQueue.scala 130:72:@11462.4]
  wire  _T_11521; // @[AxiLoadQueue.scala 131:33:@11463.4]
  wire  _T_11524; // @[AxiLoadQueue.scala 131:41:@11465.4]
  wire  _T_11526; // @[AxiLoadQueue.scala 131:9:@11466.4]
  wire  storesToCheck_15_13; // @[AxiLoadQueue.scala 130:10:@11467.4]
  wire  _T_11532; // @[AxiLoadQueue.scala 130:81:@11470.4]
  wire  _T_11533; // @[AxiLoadQueue.scala 130:72:@11471.4]
  wire  _T_11535; // @[AxiLoadQueue.scala 131:33:@11472.4]
  wire  _T_11538; // @[AxiLoadQueue.scala 131:41:@11474.4]
  wire  _T_11540; // @[AxiLoadQueue.scala 131:9:@11475.4]
  wire  storesToCheck_15_14; // @[AxiLoadQueue.scala 130:10:@11476.4]
  wire  _T_11546; // @[AxiLoadQueue.scala 130:81:@11479.4]
  wire  storesToCheck_15_15; // @[AxiLoadQueue.scala 130:10:@11485.4]
  wire  _T_12808; // @[AxiLoadQueue.scala 140:18:@11520.4]
  wire  entriesToCheck_0_0; // @[AxiLoadQueue.scala 140:26:@11521.4]
  wire  _T_12810; // @[AxiLoadQueue.scala 140:18:@11522.4]
  wire  entriesToCheck_0_1; // @[AxiLoadQueue.scala 140:26:@11523.4]
  wire  _T_12812; // @[AxiLoadQueue.scala 140:18:@11524.4]
  wire  entriesToCheck_0_2; // @[AxiLoadQueue.scala 140:26:@11525.4]
  wire  _T_12814; // @[AxiLoadQueue.scala 140:18:@11526.4]
  wire  entriesToCheck_0_3; // @[AxiLoadQueue.scala 140:26:@11527.4]
  wire  _T_12816; // @[AxiLoadQueue.scala 140:18:@11528.4]
  wire  entriesToCheck_0_4; // @[AxiLoadQueue.scala 140:26:@11529.4]
  wire  _T_12818; // @[AxiLoadQueue.scala 140:18:@11530.4]
  wire  entriesToCheck_0_5; // @[AxiLoadQueue.scala 140:26:@11531.4]
  wire  _T_12820; // @[AxiLoadQueue.scala 140:18:@11532.4]
  wire  entriesToCheck_0_6; // @[AxiLoadQueue.scala 140:26:@11533.4]
  wire  _T_12822; // @[AxiLoadQueue.scala 140:18:@11534.4]
  wire  entriesToCheck_0_7; // @[AxiLoadQueue.scala 140:26:@11535.4]
  wire  _T_12824; // @[AxiLoadQueue.scala 140:18:@11536.4]
  wire  entriesToCheck_0_8; // @[AxiLoadQueue.scala 140:26:@11537.4]
  wire  _T_12826; // @[AxiLoadQueue.scala 140:18:@11538.4]
  wire  entriesToCheck_0_9; // @[AxiLoadQueue.scala 140:26:@11539.4]
  wire  _T_12828; // @[AxiLoadQueue.scala 140:18:@11540.4]
  wire  entriesToCheck_0_10; // @[AxiLoadQueue.scala 140:26:@11541.4]
  wire  _T_12830; // @[AxiLoadQueue.scala 140:18:@11542.4]
  wire  entriesToCheck_0_11; // @[AxiLoadQueue.scala 140:26:@11543.4]
  wire  _T_12832; // @[AxiLoadQueue.scala 140:18:@11544.4]
  wire  entriesToCheck_0_12; // @[AxiLoadQueue.scala 140:26:@11545.4]
  wire  _T_12834; // @[AxiLoadQueue.scala 140:18:@11546.4]
  wire  entriesToCheck_0_13; // @[AxiLoadQueue.scala 140:26:@11547.4]
  wire  _T_12836; // @[AxiLoadQueue.scala 140:18:@11548.4]
  wire  entriesToCheck_0_14; // @[AxiLoadQueue.scala 140:26:@11549.4]
  wire  _T_12838; // @[AxiLoadQueue.scala 140:18:@11550.4]
  wire  entriesToCheck_0_15; // @[AxiLoadQueue.scala 140:26:@11551.4]
  wire  _T_12840; // @[AxiLoadQueue.scala 140:18:@11568.4]
  wire  entriesToCheck_1_0; // @[AxiLoadQueue.scala 140:26:@11569.4]
  wire  _T_12842; // @[AxiLoadQueue.scala 140:18:@11570.4]
  wire  entriesToCheck_1_1; // @[AxiLoadQueue.scala 140:26:@11571.4]
  wire  _T_12844; // @[AxiLoadQueue.scala 140:18:@11572.4]
  wire  entriesToCheck_1_2; // @[AxiLoadQueue.scala 140:26:@11573.4]
  wire  _T_12846; // @[AxiLoadQueue.scala 140:18:@11574.4]
  wire  entriesToCheck_1_3; // @[AxiLoadQueue.scala 140:26:@11575.4]
  wire  _T_12848; // @[AxiLoadQueue.scala 140:18:@11576.4]
  wire  entriesToCheck_1_4; // @[AxiLoadQueue.scala 140:26:@11577.4]
  wire  _T_12850; // @[AxiLoadQueue.scala 140:18:@11578.4]
  wire  entriesToCheck_1_5; // @[AxiLoadQueue.scala 140:26:@11579.4]
  wire  _T_12852; // @[AxiLoadQueue.scala 140:18:@11580.4]
  wire  entriesToCheck_1_6; // @[AxiLoadQueue.scala 140:26:@11581.4]
  wire  _T_12854; // @[AxiLoadQueue.scala 140:18:@11582.4]
  wire  entriesToCheck_1_7; // @[AxiLoadQueue.scala 140:26:@11583.4]
  wire  _T_12856; // @[AxiLoadQueue.scala 140:18:@11584.4]
  wire  entriesToCheck_1_8; // @[AxiLoadQueue.scala 140:26:@11585.4]
  wire  _T_12858; // @[AxiLoadQueue.scala 140:18:@11586.4]
  wire  entriesToCheck_1_9; // @[AxiLoadQueue.scala 140:26:@11587.4]
  wire  _T_12860; // @[AxiLoadQueue.scala 140:18:@11588.4]
  wire  entriesToCheck_1_10; // @[AxiLoadQueue.scala 140:26:@11589.4]
  wire  _T_12862; // @[AxiLoadQueue.scala 140:18:@11590.4]
  wire  entriesToCheck_1_11; // @[AxiLoadQueue.scala 140:26:@11591.4]
  wire  _T_12864; // @[AxiLoadQueue.scala 140:18:@11592.4]
  wire  entriesToCheck_1_12; // @[AxiLoadQueue.scala 140:26:@11593.4]
  wire  _T_12866; // @[AxiLoadQueue.scala 140:18:@11594.4]
  wire  entriesToCheck_1_13; // @[AxiLoadQueue.scala 140:26:@11595.4]
  wire  _T_12868; // @[AxiLoadQueue.scala 140:18:@11596.4]
  wire  entriesToCheck_1_14; // @[AxiLoadQueue.scala 140:26:@11597.4]
  wire  _T_12870; // @[AxiLoadQueue.scala 140:18:@11598.4]
  wire  entriesToCheck_1_15; // @[AxiLoadQueue.scala 140:26:@11599.4]
  wire  _T_12872; // @[AxiLoadQueue.scala 140:18:@11616.4]
  wire  entriesToCheck_2_0; // @[AxiLoadQueue.scala 140:26:@11617.4]
  wire  _T_12874; // @[AxiLoadQueue.scala 140:18:@11618.4]
  wire  entriesToCheck_2_1; // @[AxiLoadQueue.scala 140:26:@11619.4]
  wire  _T_12876; // @[AxiLoadQueue.scala 140:18:@11620.4]
  wire  entriesToCheck_2_2; // @[AxiLoadQueue.scala 140:26:@11621.4]
  wire  _T_12878; // @[AxiLoadQueue.scala 140:18:@11622.4]
  wire  entriesToCheck_2_3; // @[AxiLoadQueue.scala 140:26:@11623.4]
  wire  _T_12880; // @[AxiLoadQueue.scala 140:18:@11624.4]
  wire  entriesToCheck_2_4; // @[AxiLoadQueue.scala 140:26:@11625.4]
  wire  _T_12882; // @[AxiLoadQueue.scala 140:18:@11626.4]
  wire  entriesToCheck_2_5; // @[AxiLoadQueue.scala 140:26:@11627.4]
  wire  _T_12884; // @[AxiLoadQueue.scala 140:18:@11628.4]
  wire  entriesToCheck_2_6; // @[AxiLoadQueue.scala 140:26:@11629.4]
  wire  _T_12886; // @[AxiLoadQueue.scala 140:18:@11630.4]
  wire  entriesToCheck_2_7; // @[AxiLoadQueue.scala 140:26:@11631.4]
  wire  _T_12888; // @[AxiLoadQueue.scala 140:18:@11632.4]
  wire  entriesToCheck_2_8; // @[AxiLoadQueue.scala 140:26:@11633.4]
  wire  _T_12890; // @[AxiLoadQueue.scala 140:18:@11634.4]
  wire  entriesToCheck_2_9; // @[AxiLoadQueue.scala 140:26:@11635.4]
  wire  _T_12892; // @[AxiLoadQueue.scala 140:18:@11636.4]
  wire  entriesToCheck_2_10; // @[AxiLoadQueue.scala 140:26:@11637.4]
  wire  _T_12894; // @[AxiLoadQueue.scala 140:18:@11638.4]
  wire  entriesToCheck_2_11; // @[AxiLoadQueue.scala 140:26:@11639.4]
  wire  _T_12896; // @[AxiLoadQueue.scala 140:18:@11640.4]
  wire  entriesToCheck_2_12; // @[AxiLoadQueue.scala 140:26:@11641.4]
  wire  _T_12898; // @[AxiLoadQueue.scala 140:18:@11642.4]
  wire  entriesToCheck_2_13; // @[AxiLoadQueue.scala 140:26:@11643.4]
  wire  _T_12900; // @[AxiLoadQueue.scala 140:18:@11644.4]
  wire  entriesToCheck_2_14; // @[AxiLoadQueue.scala 140:26:@11645.4]
  wire  _T_12902; // @[AxiLoadQueue.scala 140:18:@11646.4]
  wire  entriesToCheck_2_15; // @[AxiLoadQueue.scala 140:26:@11647.4]
  wire  _T_12904; // @[AxiLoadQueue.scala 140:18:@11664.4]
  wire  entriesToCheck_3_0; // @[AxiLoadQueue.scala 140:26:@11665.4]
  wire  _T_12906; // @[AxiLoadQueue.scala 140:18:@11666.4]
  wire  entriesToCheck_3_1; // @[AxiLoadQueue.scala 140:26:@11667.4]
  wire  _T_12908; // @[AxiLoadQueue.scala 140:18:@11668.4]
  wire  entriesToCheck_3_2; // @[AxiLoadQueue.scala 140:26:@11669.4]
  wire  _T_12910; // @[AxiLoadQueue.scala 140:18:@11670.4]
  wire  entriesToCheck_3_3; // @[AxiLoadQueue.scala 140:26:@11671.4]
  wire  _T_12912; // @[AxiLoadQueue.scala 140:18:@11672.4]
  wire  entriesToCheck_3_4; // @[AxiLoadQueue.scala 140:26:@11673.4]
  wire  _T_12914; // @[AxiLoadQueue.scala 140:18:@11674.4]
  wire  entriesToCheck_3_5; // @[AxiLoadQueue.scala 140:26:@11675.4]
  wire  _T_12916; // @[AxiLoadQueue.scala 140:18:@11676.4]
  wire  entriesToCheck_3_6; // @[AxiLoadQueue.scala 140:26:@11677.4]
  wire  _T_12918; // @[AxiLoadQueue.scala 140:18:@11678.4]
  wire  entriesToCheck_3_7; // @[AxiLoadQueue.scala 140:26:@11679.4]
  wire  _T_12920; // @[AxiLoadQueue.scala 140:18:@11680.4]
  wire  entriesToCheck_3_8; // @[AxiLoadQueue.scala 140:26:@11681.4]
  wire  _T_12922; // @[AxiLoadQueue.scala 140:18:@11682.4]
  wire  entriesToCheck_3_9; // @[AxiLoadQueue.scala 140:26:@11683.4]
  wire  _T_12924; // @[AxiLoadQueue.scala 140:18:@11684.4]
  wire  entriesToCheck_3_10; // @[AxiLoadQueue.scala 140:26:@11685.4]
  wire  _T_12926; // @[AxiLoadQueue.scala 140:18:@11686.4]
  wire  entriesToCheck_3_11; // @[AxiLoadQueue.scala 140:26:@11687.4]
  wire  _T_12928; // @[AxiLoadQueue.scala 140:18:@11688.4]
  wire  entriesToCheck_3_12; // @[AxiLoadQueue.scala 140:26:@11689.4]
  wire  _T_12930; // @[AxiLoadQueue.scala 140:18:@11690.4]
  wire  entriesToCheck_3_13; // @[AxiLoadQueue.scala 140:26:@11691.4]
  wire  _T_12932; // @[AxiLoadQueue.scala 140:18:@11692.4]
  wire  entriesToCheck_3_14; // @[AxiLoadQueue.scala 140:26:@11693.4]
  wire  _T_12934; // @[AxiLoadQueue.scala 140:18:@11694.4]
  wire  entriesToCheck_3_15; // @[AxiLoadQueue.scala 140:26:@11695.4]
  wire  _T_12936; // @[AxiLoadQueue.scala 140:18:@11712.4]
  wire  entriesToCheck_4_0; // @[AxiLoadQueue.scala 140:26:@11713.4]
  wire  _T_12938; // @[AxiLoadQueue.scala 140:18:@11714.4]
  wire  entriesToCheck_4_1; // @[AxiLoadQueue.scala 140:26:@11715.4]
  wire  _T_12940; // @[AxiLoadQueue.scala 140:18:@11716.4]
  wire  entriesToCheck_4_2; // @[AxiLoadQueue.scala 140:26:@11717.4]
  wire  _T_12942; // @[AxiLoadQueue.scala 140:18:@11718.4]
  wire  entriesToCheck_4_3; // @[AxiLoadQueue.scala 140:26:@11719.4]
  wire  _T_12944; // @[AxiLoadQueue.scala 140:18:@11720.4]
  wire  entriesToCheck_4_4; // @[AxiLoadQueue.scala 140:26:@11721.4]
  wire  _T_12946; // @[AxiLoadQueue.scala 140:18:@11722.4]
  wire  entriesToCheck_4_5; // @[AxiLoadQueue.scala 140:26:@11723.4]
  wire  _T_12948; // @[AxiLoadQueue.scala 140:18:@11724.4]
  wire  entriesToCheck_4_6; // @[AxiLoadQueue.scala 140:26:@11725.4]
  wire  _T_12950; // @[AxiLoadQueue.scala 140:18:@11726.4]
  wire  entriesToCheck_4_7; // @[AxiLoadQueue.scala 140:26:@11727.4]
  wire  _T_12952; // @[AxiLoadQueue.scala 140:18:@11728.4]
  wire  entriesToCheck_4_8; // @[AxiLoadQueue.scala 140:26:@11729.4]
  wire  _T_12954; // @[AxiLoadQueue.scala 140:18:@11730.4]
  wire  entriesToCheck_4_9; // @[AxiLoadQueue.scala 140:26:@11731.4]
  wire  _T_12956; // @[AxiLoadQueue.scala 140:18:@11732.4]
  wire  entriesToCheck_4_10; // @[AxiLoadQueue.scala 140:26:@11733.4]
  wire  _T_12958; // @[AxiLoadQueue.scala 140:18:@11734.4]
  wire  entriesToCheck_4_11; // @[AxiLoadQueue.scala 140:26:@11735.4]
  wire  _T_12960; // @[AxiLoadQueue.scala 140:18:@11736.4]
  wire  entriesToCheck_4_12; // @[AxiLoadQueue.scala 140:26:@11737.4]
  wire  _T_12962; // @[AxiLoadQueue.scala 140:18:@11738.4]
  wire  entriesToCheck_4_13; // @[AxiLoadQueue.scala 140:26:@11739.4]
  wire  _T_12964; // @[AxiLoadQueue.scala 140:18:@11740.4]
  wire  entriesToCheck_4_14; // @[AxiLoadQueue.scala 140:26:@11741.4]
  wire  _T_12966; // @[AxiLoadQueue.scala 140:18:@11742.4]
  wire  entriesToCheck_4_15; // @[AxiLoadQueue.scala 140:26:@11743.4]
  wire  _T_12968; // @[AxiLoadQueue.scala 140:18:@11760.4]
  wire  entriesToCheck_5_0; // @[AxiLoadQueue.scala 140:26:@11761.4]
  wire  _T_12970; // @[AxiLoadQueue.scala 140:18:@11762.4]
  wire  entriesToCheck_5_1; // @[AxiLoadQueue.scala 140:26:@11763.4]
  wire  _T_12972; // @[AxiLoadQueue.scala 140:18:@11764.4]
  wire  entriesToCheck_5_2; // @[AxiLoadQueue.scala 140:26:@11765.4]
  wire  _T_12974; // @[AxiLoadQueue.scala 140:18:@11766.4]
  wire  entriesToCheck_5_3; // @[AxiLoadQueue.scala 140:26:@11767.4]
  wire  _T_12976; // @[AxiLoadQueue.scala 140:18:@11768.4]
  wire  entriesToCheck_5_4; // @[AxiLoadQueue.scala 140:26:@11769.4]
  wire  _T_12978; // @[AxiLoadQueue.scala 140:18:@11770.4]
  wire  entriesToCheck_5_5; // @[AxiLoadQueue.scala 140:26:@11771.4]
  wire  _T_12980; // @[AxiLoadQueue.scala 140:18:@11772.4]
  wire  entriesToCheck_5_6; // @[AxiLoadQueue.scala 140:26:@11773.4]
  wire  _T_12982; // @[AxiLoadQueue.scala 140:18:@11774.4]
  wire  entriesToCheck_5_7; // @[AxiLoadQueue.scala 140:26:@11775.4]
  wire  _T_12984; // @[AxiLoadQueue.scala 140:18:@11776.4]
  wire  entriesToCheck_5_8; // @[AxiLoadQueue.scala 140:26:@11777.4]
  wire  _T_12986; // @[AxiLoadQueue.scala 140:18:@11778.4]
  wire  entriesToCheck_5_9; // @[AxiLoadQueue.scala 140:26:@11779.4]
  wire  _T_12988; // @[AxiLoadQueue.scala 140:18:@11780.4]
  wire  entriesToCheck_5_10; // @[AxiLoadQueue.scala 140:26:@11781.4]
  wire  _T_12990; // @[AxiLoadQueue.scala 140:18:@11782.4]
  wire  entriesToCheck_5_11; // @[AxiLoadQueue.scala 140:26:@11783.4]
  wire  _T_12992; // @[AxiLoadQueue.scala 140:18:@11784.4]
  wire  entriesToCheck_5_12; // @[AxiLoadQueue.scala 140:26:@11785.4]
  wire  _T_12994; // @[AxiLoadQueue.scala 140:18:@11786.4]
  wire  entriesToCheck_5_13; // @[AxiLoadQueue.scala 140:26:@11787.4]
  wire  _T_12996; // @[AxiLoadQueue.scala 140:18:@11788.4]
  wire  entriesToCheck_5_14; // @[AxiLoadQueue.scala 140:26:@11789.4]
  wire  _T_12998; // @[AxiLoadQueue.scala 140:18:@11790.4]
  wire  entriesToCheck_5_15; // @[AxiLoadQueue.scala 140:26:@11791.4]
  wire  _T_13000; // @[AxiLoadQueue.scala 140:18:@11808.4]
  wire  entriesToCheck_6_0; // @[AxiLoadQueue.scala 140:26:@11809.4]
  wire  _T_13002; // @[AxiLoadQueue.scala 140:18:@11810.4]
  wire  entriesToCheck_6_1; // @[AxiLoadQueue.scala 140:26:@11811.4]
  wire  _T_13004; // @[AxiLoadQueue.scala 140:18:@11812.4]
  wire  entriesToCheck_6_2; // @[AxiLoadQueue.scala 140:26:@11813.4]
  wire  _T_13006; // @[AxiLoadQueue.scala 140:18:@11814.4]
  wire  entriesToCheck_6_3; // @[AxiLoadQueue.scala 140:26:@11815.4]
  wire  _T_13008; // @[AxiLoadQueue.scala 140:18:@11816.4]
  wire  entriesToCheck_6_4; // @[AxiLoadQueue.scala 140:26:@11817.4]
  wire  _T_13010; // @[AxiLoadQueue.scala 140:18:@11818.4]
  wire  entriesToCheck_6_5; // @[AxiLoadQueue.scala 140:26:@11819.4]
  wire  _T_13012; // @[AxiLoadQueue.scala 140:18:@11820.4]
  wire  entriesToCheck_6_6; // @[AxiLoadQueue.scala 140:26:@11821.4]
  wire  _T_13014; // @[AxiLoadQueue.scala 140:18:@11822.4]
  wire  entriesToCheck_6_7; // @[AxiLoadQueue.scala 140:26:@11823.4]
  wire  _T_13016; // @[AxiLoadQueue.scala 140:18:@11824.4]
  wire  entriesToCheck_6_8; // @[AxiLoadQueue.scala 140:26:@11825.4]
  wire  _T_13018; // @[AxiLoadQueue.scala 140:18:@11826.4]
  wire  entriesToCheck_6_9; // @[AxiLoadQueue.scala 140:26:@11827.4]
  wire  _T_13020; // @[AxiLoadQueue.scala 140:18:@11828.4]
  wire  entriesToCheck_6_10; // @[AxiLoadQueue.scala 140:26:@11829.4]
  wire  _T_13022; // @[AxiLoadQueue.scala 140:18:@11830.4]
  wire  entriesToCheck_6_11; // @[AxiLoadQueue.scala 140:26:@11831.4]
  wire  _T_13024; // @[AxiLoadQueue.scala 140:18:@11832.4]
  wire  entriesToCheck_6_12; // @[AxiLoadQueue.scala 140:26:@11833.4]
  wire  _T_13026; // @[AxiLoadQueue.scala 140:18:@11834.4]
  wire  entriesToCheck_6_13; // @[AxiLoadQueue.scala 140:26:@11835.4]
  wire  _T_13028; // @[AxiLoadQueue.scala 140:18:@11836.4]
  wire  entriesToCheck_6_14; // @[AxiLoadQueue.scala 140:26:@11837.4]
  wire  _T_13030; // @[AxiLoadQueue.scala 140:18:@11838.4]
  wire  entriesToCheck_6_15; // @[AxiLoadQueue.scala 140:26:@11839.4]
  wire  _T_13032; // @[AxiLoadQueue.scala 140:18:@11856.4]
  wire  entriesToCheck_7_0; // @[AxiLoadQueue.scala 140:26:@11857.4]
  wire  _T_13034; // @[AxiLoadQueue.scala 140:18:@11858.4]
  wire  entriesToCheck_7_1; // @[AxiLoadQueue.scala 140:26:@11859.4]
  wire  _T_13036; // @[AxiLoadQueue.scala 140:18:@11860.4]
  wire  entriesToCheck_7_2; // @[AxiLoadQueue.scala 140:26:@11861.4]
  wire  _T_13038; // @[AxiLoadQueue.scala 140:18:@11862.4]
  wire  entriesToCheck_7_3; // @[AxiLoadQueue.scala 140:26:@11863.4]
  wire  _T_13040; // @[AxiLoadQueue.scala 140:18:@11864.4]
  wire  entriesToCheck_7_4; // @[AxiLoadQueue.scala 140:26:@11865.4]
  wire  _T_13042; // @[AxiLoadQueue.scala 140:18:@11866.4]
  wire  entriesToCheck_7_5; // @[AxiLoadQueue.scala 140:26:@11867.4]
  wire  _T_13044; // @[AxiLoadQueue.scala 140:18:@11868.4]
  wire  entriesToCheck_7_6; // @[AxiLoadQueue.scala 140:26:@11869.4]
  wire  _T_13046; // @[AxiLoadQueue.scala 140:18:@11870.4]
  wire  entriesToCheck_7_7; // @[AxiLoadQueue.scala 140:26:@11871.4]
  wire  _T_13048; // @[AxiLoadQueue.scala 140:18:@11872.4]
  wire  entriesToCheck_7_8; // @[AxiLoadQueue.scala 140:26:@11873.4]
  wire  _T_13050; // @[AxiLoadQueue.scala 140:18:@11874.4]
  wire  entriesToCheck_7_9; // @[AxiLoadQueue.scala 140:26:@11875.4]
  wire  _T_13052; // @[AxiLoadQueue.scala 140:18:@11876.4]
  wire  entriesToCheck_7_10; // @[AxiLoadQueue.scala 140:26:@11877.4]
  wire  _T_13054; // @[AxiLoadQueue.scala 140:18:@11878.4]
  wire  entriesToCheck_7_11; // @[AxiLoadQueue.scala 140:26:@11879.4]
  wire  _T_13056; // @[AxiLoadQueue.scala 140:18:@11880.4]
  wire  entriesToCheck_7_12; // @[AxiLoadQueue.scala 140:26:@11881.4]
  wire  _T_13058; // @[AxiLoadQueue.scala 140:18:@11882.4]
  wire  entriesToCheck_7_13; // @[AxiLoadQueue.scala 140:26:@11883.4]
  wire  _T_13060; // @[AxiLoadQueue.scala 140:18:@11884.4]
  wire  entriesToCheck_7_14; // @[AxiLoadQueue.scala 140:26:@11885.4]
  wire  _T_13062; // @[AxiLoadQueue.scala 140:18:@11886.4]
  wire  entriesToCheck_7_15; // @[AxiLoadQueue.scala 140:26:@11887.4]
  wire  _T_13064; // @[AxiLoadQueue.scala 140:18:@11904.4]
  wire  entriesToCheck_8_0; // @[AxiLoadQueue.scala 140:26:@11905.4]
  wire  _T_13066; // @[AxiLoadQueue.scala 140:18:@11906.4]
  wire  entriesToCheck_8_1; // @[AxiLoadQueue.scala 140:26:@11907.4]
  wire  _T_13068; // @[AxiLoadQueue.scala 140:18:@11908.4]
  wire  entriesToCheck_8_2; // @[AxiLoadQueue.scala 140:26:@11909.4]
  wire  _T_13070; // @[AxiLoadQueue.scala 140:18:@11910.4]
  wire  entriesToCheck_8_3; // @[AxiLoadQueue.scala 140:26:@11911.4]
  wire  _T_13072; // @[AxiLoadQueue.scala 140:18:@11912.4]
  wire  entriesToCheck_8_4; // @[AxiLoadQueue.scala 140:26:@11913.4]
  wire  _T_13074; // @[AxiLoadQueue.scala 140:18:@11914.4]
  wire  entriesToCheck_8_5; // @[AxiLoadQueue.scala 140:26:@11915.4]
  wire  _T_13076; // @[AxiLoadQueue.scala 140:18:@11916.4]
  wire  entriesToCheck_8_6; // @[AxiLoadQueue.scala 140:26:@11917.4]
  wire  _T_13078; // @[AxiLoadQueue.scala 140:18:@11918.4]
  wire  entriesToCheck_8_7; // @[AxiLoadQueue.scala 140:26:@11919.4]
  wire  _T_13080; // @[AxiLoadQueue.scala 140:18:@11920.4]
  wire  entriesToCheck_8_8; // @[AxiLoadQueue.scala 140:26:@11921.4]
  wire  _T_13082; // @[AxiLoadQueue.scala 140:18:@11922.4]
  wire  entriesToCheck_8_9; // @[AxiLoadQueue.scala 140:26:@11923.4]
  wire  _T_13084; // @[AxiLoadQueue.scala 140:18:@11924.4]
  wire  entriesToCheck_8_10; // @[AxiLoadQueue.scala 140:26:@11925.4]
  wire  _T_13086; // @[AxiLoadQueue.scala 140:18:@11926.4]
  wire  entriesToCheck_8_11; // @[AxiLoadQueue.scala 140:26:@11927.4]
  wire  _T_13088; // @[AxiLoadQueue.scala 140:18:@11928.4]
  wire  entriesToCheck_8_12; // @[AxiLoadQueue.scala 140:26:@11929.4]
  wire  _T_13090; // @[AxiLoadQueue.scala 140:18:@11930.4]
  wire  entriesToCheck_8_13; // @[AxiLoadQueue.scala 140:26:@11931.4]
  wire  _T_13092; // @[AxiLoadQueue.scala 140:18:@11932.4]
  wire  entriesToCheck_8_14; // @[AxiLoadQueue.scala 140:26:@11933.4]
  wire  _T_13094; // @[AxiLoadQueue.scala 140:18:@11934.4]
  wire  entriesToCheck_8_15; // @[AxiLoadQueue.scala 140:26:@11935.4]
  wire  _T_13096; // @[AxiLoadQueue.scala 140:18:@11952.4]
  wire  entriesToCheck_9_0; // @[AxiLoadQueue.scala 140:26:@11953.4]
  wire  _T_13098; // @[AxiLoadQueue.scala 140:18:@11954.4]
  wire  entriesToCheck_9_1; // @[AxiLoadQueue.scala 140:26:@11955.4]
  wire  _T_13100; // @[AxiLoadQueue.scala 140:18:@11956.4]
  wire  entriesToCheck_9_2; // @[AxiLoadQueue.scala 140:26:@11957.4]
  wire  _T_13102; // @[AxiLoadQueue.scala 140:18:@11958.4]
  wire  entriesToCheck_9_3; // @[AxiLoadQueue.scala 140:26:@11959.4]
  wire  _T_13104; // @[AxiLoadQueue.scala 140:18:@11960.4]
  wire  entriesToCheck_9_4; // @[AxiLoadQueue.scala 140:26:@11961.4]
  wire  _T_13106; // @[AxiLoadQueue.scala 140:18:@11962.4]
  wire  entriesToCheck_9_5; // @[AxiLoadQueue.scala 140:26:@11963.4]
  wire  _T_13108; // @[AxiLoadQueue.scala 140:18:@11964.4]
  wire  entriesToCheck_9_6; // @[AxiLoadQueue.scala 140:26:@11965.4]
  wire  _T_13110; // @[AxiLoadQueue.scala 140:18:@11966.4]
  wire  entriesToCheck_9_7; // @[AxiLoadQueue.scala 140:26:@11967.4]
  wire  _T_13112; // @[AxiLoadQueue.scala 140:18:@11968.4]
  wire  entriesToCheck_9_8; // @[AxiLoadQueue.scala 140:26:@11969.4]
  wire  _T_13114; // @[AxiLoadQueue.scala 140:18:@11970.4]
  wire  entriesToCheck_9_9; // @[AxiLoadQueue.scala 140:26:@11971.4]
  wire  _T_13116; // @[AxiLoadQueue.scala 140:18:@11972.4]
  wire  entriesToCheck_9_10; // @[AxiLoadQueue.scala 140:26:@11973.4]
  wire  _T_13118; // @[AxiLoadQueue.scala 140:18:@11974.4]
  wire  entriesToCheck_9_11; // @[AxiLoadQueue.scala 140:26:@11975.4]
  wire  _T_13120; // @[AxiLoadQueue.scala 140:18:@11976.4]
  wire  entriesToCheck_9_12; // @[AxiLoadQueue.scala 140:26:@11977.4]
  wire  _T_13122; // @[AxiLoadQueue.scala 140:18:@11978.4]
  wire  entriesToCheck_9_13; // @[AxiLoadQueue.scala 140:26:@11979.4]
  wire  _T_13124; // @[AxiLoadQueue.scala 140:18:@11980.4]
  wire  entriesToCheck_9_14; // @[AxiLoadQueue.scala 140:26:@11981.4]
  wire  _T_13126; // @[AxiLoadQueue.scala 140:18:@11982.4]
  wire  entriesToCheck_9_15; // @[AxiLoadQueue.scala 140:26:@11983.4]
  wire  _T_13128; // @[AxiLoadQueue.scala 140:18:@12000.4]
  wire  entriesToCheck_10_0; // @[AxiLoadQueue.scala 140:26:@12001.4]
  wire  _T_13130; // @[AxiLoadQueue.scala 140:18:@12002.4]
  wire  entriesToCheck_10_1; // @[AxiLoadQueue.scala 140:26:@12003.4]
  wire  _T_13132; // @[AxiLoadQueue.scala 140:18:@12004.4]
  wire  entriesToCheck_10_2; // @[AxiLoadQueue.scala 140:26:@12005.4]
  wire  _T_13134; // @[AxiLoadQueue.scala 140:18:@12006.4]
  wire  entriesToCheck_10_3; // @[AxiLoadQueue.scala 140:26:@12007.4]
  wire  _T_13136; // @[AxiLoadQueue.scala 140:18:@12008.4]
  wire  entriesToCheck_10_4; // @[AxiLoadQueue.scala 140:26:@12009.4]
  wire  _T_13138; // @[AxiLoadQueue.scala 140:18:@12010.4]
  wire  entriesToCheck_10_5; // @[AxiLoadQueue.scala 140:26:@12011.4]
  wire  _T_13140; // @[AxiLoadQueue.scala 140:18:@12012.4]
  wire  entriesToCheck_10_6; // @[AxiLoadQueue.scala 140:26:@12013.4]
  wire  _T_13142; // @[AxiLoadQueue.scala 140:18:@12014.4]
  wire  entriesToCheck_10_7; // @[AxiLoadQueue.scala 140:26:@12015.4]
  wire  _T_13144; // @[AxiLoadQueue.scala 140:18:@12016.4]
  wire  entriesToCheck_10_8; // @[AxiLoadQueue.scala 140:26:@12017.4]
  wire  _T_13146; // @[AxiLoadQueue.scala 140:18:@12018.4]
  wire  entriesToCheck_10_9; // @[AxiLoadQueue.scala 140:26:@12019.4]
  wire  _T_13148; // @[AxiLoadQueue.scala 140:18:@12020.4]
  wire  entriesToCheck_10_10; // @[AxiLoadQueue.scala 140:26:@12021.4]
  wire  _T_13150; // @[AxiLoadQueue.scala 140:18:@12022.4]
  wire  entriesToCheck_10_11; // @[AxiLoadQueue.scala 140:26:@12023.4]
  wire  _T_13152; // @[AxiLoadQueue.scala 140:18:@12024.4]
  wire  entriesToCheck_10_12; // @[AxiLoadQueue.scala 140:26:@12025.4]
  wire  _T_13154; // @[AxiLoadQueue.scala 140:18:@12026.4]
  wire  entriesToCheck_10_13; // @[AxiLoadQueue.scala 140:26:@12027.4]
  wire  _T_13156; // @[AxiLoadQueue.scala 140:18:@12028.4]
  wire  entriesToCheck_10_14; // @[AxiLoadQueue.scala 140:26:@12029.4]
  wire  _T_13158; // @[AxiLoadQueue.scala 140:18:@12030.4]
  wire  entriesToCheck_10_15; // @[AxiLoadQueue.scala 140:26:@12031.4]
  wire  _T_13160; // @[AxiLoadQueue.scala 140:18:@12048.4]
  wire  entriesToCheck_11_0; // @[AxiLoadQueue.scala 140:26:@12049.4]
  wire  _T_13162; // @[AxiLoadQueue.scala 140:18:@12050.4]
  wire  entriesToCheck_11_1; // @[AxiLoadQueue.scala 140:26:@12051.4]
  wire  _T_13164; // @[AxiLoadQueue.scala 140:18:@12052.4]
  wire  entriesToCheck_11_2; // @[AxiLoadQueue.scala 140:26:@12053.4]
  wire  _T_13166; // @[AxiLoadQueue.scala 140:18:@12054.4]
  wire  entriesToCheck_11_3; // @[AxiLoadQueue.scala 140:26:@12055.4]
  wire  _T_13168; // @[AxiLoadQueue.scala 140:18:@12056.4]
  wire  entriesToCheck_11_4; // @[AxiLoadQueue.scala 140:26:@12057.4]
  wire  _T_13170; // @[AxiLoadQueue.scala 140:18:@12058.4]
  wire  entriesToCheck_11_5; // @[AxiLoadQueue.scala 140:26:@12059.4]
  wire  _T_13172; // @[AxiLoadQueue.scala 140:18:@12060.4]
  wire  entriesToCheck_11_6; // @[AxiLoadQueue.scala 140:26:@12061.4]
  wire  _T_13174; // @[AxiLoadQueue.scala 140:18:@12062.4]
  wire  entriesToCheck_11_7; // @[AxiLoadQueue.scala 140:26:@12063.4]
  wire  _T_13176; // @[AxiLoadQueue.scala 140:18:@12064.4]
  wire  entriesToCheck_11_8; // @[AxiLoadQueue.scala 140:26:@12065.4]
  wire  _T_13178; // @[AxiLoadQueue.scala 140:18:@12066.4]
  wire  entriesToCheck_11_9; // @[AxiLoadQueue.scala 140:26:@12067.4]
  wire  _T_13180; // @[AxiLoadQueue.scala 140:18:@12068.4]
  wire  entriesToCheck_11_10; // @[AxiLoadQueue.scala 140:26:@12069.4]
  wire  _T_13182; // @[AxiLoadQueue.scala 140:18:@12070.4]
  wire  entriesToCheck_11_11; // @[AxiLoadQueue.scala 140:26:@12071.4]
  wire  _T_13184; // @[AxiLoadQueue.scala 140:18:@12072.4]
  wire  entriesToCheck_11_12; // @[AxiLoadQueue.scala 140:26:@12073.4]
  wire  _T_13186; // @[AxiLoadQueue.scala 140:18:@12074.4]
  wire  entriesToCheck_11_13; // @[AxiLoadQueue.scala 140:26:@12075.4]
  wire  _T_13188; // @[AxiLoadQueue.scala 140:18:@12076.4]
  wire  entriesToCheck_11_14; // @[AxiLoadQueue.scala 140:26:@12077.4]
  wire  _T_13190; // @[AxiLoadQueue.scala 140:18:@12078.4]
  wire  entriesToCheck_11_15; // @[AxiLoadQueue.scala 140:26:@12079.4]
  wire  _T_13192; // @[AxiLoadQueue.scala 140:18:@12096.4]
  wire  entriesToCheck_12_0; // @[AxiLoadQueue.scala 140:26:@12097.4]
  wire  _T_13194; // @[AxiLoadQueue.scala 140:18:@12098.4]
  wire  entriesToCheck_12_1; // @[AxiLoadQueue.scala 140:26:@12099.4]
  wire  _T_13196; // @[AxiLoadQueue.scala 140:18:@12100.4]
  wire  entriesToCheck_12_2; // @[AxiLoadQueue.scala 140:26:@12101.4]
  wire  _T_13198; // @[AxiLoadQueue.scala 140:18:@12102.4]
  wire  entriesToCheck_12_3; // @[AxiLoadQueue.scala 140:26:@12103.4]
  wire  _T_13200; // @[AxiLoadQueue.scala 140:18:@12104.4]
  wire  entriesToCheck_12_4; // @[AxiLoadQueue.scala 140:26:@12105.4]
  wire  _T_13202; // @[AxiLoadQueue.scala 140:18:@12106.4]
  wire  entriesToCheck_12_5; // @[AxiLoadQueue.scala 140:26:@12107.4]
  wire  _T_13204; // @[AxiLoadQueue.scala 140:18:@12108.4]
  wire  entriesToCheck_12_6; // @[AxiLoadQueue.scala 140:26:@12109.4]
  wire  _T_13206; // @[AxiLoadQueue.scala 140:18:@12110.4]
  wire  entriesToCheck_12_7; // @[AxiLoadQueue.scala 140:26:@12111.4]
  wire  _T_13208; // @[AxiLoadQueue.scala 140:18:@12112.4]
  wire  entriesToCheck_12_8; // @[AxiLoadQueue.scala 140:26:@12113.4]
  wire  _T_13210; // @[AxiLoadQueue.scala 140:18:@12114.4]
  wire  entriesToCheck_12_9; // @[AxiLoadQueue.scala 140:26:@12115.4]
  wire  _T_13212; // @[AxiLoadQueue.scala 140:18:@12116.4]
  wire  entriesToCheck_12_10; // @[AxiLoadQueue.scala 140:26:@12117.4]
  wire  _T_13214; // @[AxiLoadQueue.scala 140:18:@12118.4]
  wire  entriesToCheck_12_11; // @[AxiLoadQueue.scala 140:26:@12119.4]
  wire  _T_13216; // @[AxiLoadQueue.scala 140:18:@12120.4]
  wire  entriesToCheck_12_12; // @[AxiLoadQueue.scala 140:26:@12121.4]
  wire  _T_13218; // @[AxiLoadQueue.scala 140:18:@12122.4]
  wire  entriesToCheck_12_13; // @[AxiLoadQueue.scala 140:26:@12123.4]
  wire  _T_13220; // @[AxiLoadQueue.scala 140:18:@12124.4]
  wire  entriesToCheck_12_14; // @[AxiLoadQueue.scala 140:26:@12125.4]
  wire  _T_13222; // @[AxiLoadQueue.scala 140:18:@12126.4]
  wire  entriesToCheck_12_15; // @[AxiLoadQueue.scala 140:26:@12127.4]
  wire  _T_13224; // @[AxiLoadQueue.scala 140:18:@12144.4]
  wire  entriesToCheck_13_0; // @[AxiLoadQueue.scala 140:26:@12145.4]
  wire  _T_13226; // @[AxiLoadQueue.scala 140:18:@12146.4]
  wire  entriesToCheck_13_1; // @[AxiLoadQueue.scala 140:26:@12147.4]
  wire  _T_13228; // @[AxiLoadQueue.scala 140:18:@12148.4]
  wire  entriesToCheck_13_2; // @[AxiLoadQueue.scala 140:26:@12149.4]
  wire  _T_13230; // @[AxiLoadQueue.scala 140:18:@12150.4]
  wire  entriesToCheck_13_3; // @[AxiLoadQueue.scala 140:26:@12151.4]
  wire  _T_13232; // @[AxiLoadQueue.scala 140:18:@12152.4]
  wire  entriesToCheck_13_4; // @[AxiLoadQueue.scala 140:26:@12153.4]
  wire  _T_13234; // @[AxiLoadQueue.scala 140:18:@12154.4]
  wire  entriesToCheck_13_5; // @[AxiLoadQueue.scala 140:26:@12155.4]
  wire  _T_13236; // @[AxiLoadQueue.scala 140:18:@12156.4]
  wire  entriesToCheck_13_6; // @[AxiLoadQueue.scala 140:26:@12157.4]
  wire  _T_13238; // @[AxiLoadQueue.scala 140:18:@12158.4]
  wire  entriesToCheck_13_7; // @[AxiLoadQueue.scala 140:26:@12159.4]
  wire  _T_13240; // @[AxiLoadQueue.scala 140:18:@12160.4]
  wire  entriesToCheck_13_8; // @[AxiLoadQueue.scala 140:26:@12161.4]
  wire  _T_13242; // @[AxiLoadQueue.scala 140:18:@12162.4]
  wire  entriesToCheck_13_9; // @[AxiLoadQueue.scala 140:26:@12163.4]
  wire  _T_13244; // @[AxiLoadQueue.scala 140:18:@12164.4]
  wire  entriesToCheck_13_10; // @[AxiLoadQueue.scala 140:26:@12165.4]
  wire  _T_13246; // @[AxiLoadQueue.scala 140:18:@12166.4]
  wire  entriesToCheck_13_11; // @[AxiLoadQueue.scala 140:26:@12167.4]
  wire  _T_13248; // @[AxiLoadQueue.scala 140:18:@12168.4]
  wire  entriesToCheck_13_12; // @[AxiLoadQueue.scala 140:26:@12169.4]
  wire  _T_13250; // @[AxiLoadQueue.scala 140:18:@12170.4]
  wire  entriesToCheck_13_13; // @[AxiLoadQueue.scala 140:26:@12171.4]
  wire  _T_13252; // @[AxiLoadQueue.scala 140:18:@12172.4]
  wire  entriesToCheck_13_14; // @[AxiLoadQueue.scala 140:26:@12173.4]
  wire  _T_13254; // @[AxiLoadQueue.scala 140:18:@12174.4]
  wire  entriesToCheck_13_15; // @[AxiLoadQueue.scala 140:26:@12175.4]
  wire  _T_13256; // @[AxiLoadQueue.scala 140:18:@12192.4]
  wire  entriesToCheck_14_0; // @[AxiLoadQueue.scala 140:26:@12193.4]
  wire  _T_13258; // @[AxiLoadQueue.scala 140:18:@12194.4]
  wire  entriesToCheck_14_1; // @[AxiLoadQueue.scala 140:26:@12195.4]
  wire  _T_13260; // @[AxiLoadQueue.scala 140:18:@12196.4]
  wire  entriesToCheck_14_2; // @[AxiLoadQueue.scala 140:26:@12197.4]
  wire  _T_13262; // @[AxiLoadQueue.scala 140:18:@12198.4]
  wire  entriesToCheck_14_3; // @[AxiLoadQueue.scala 140:26:@12199.4]
  wire  _T_13264; // @[AxiLoadQueue.scala 140:18:@12200.4]
  wire  entriesToCheck_14_4; // @[AxiLoadQueue.scala 140:26:@12201.4]
  wire  _T_13266; // @[AxiLoadQueue.scala 140:18:@12202.4]
  wire  entriesToCheck_14_5; // @[AxiLoadQueue.scala 140:26:@12203.4]
  wire  _T_13268; // @[AxiLoadQueue.scala 140:18:@12204.4]
  wire  entriesToCheck_14_6; // @[AxiLoadQueue.scala 140:26:@12205.4]
  wire  _T_13270; // @[AxiLoadQueue.scala 140:18:@12206.4]
  wire  entriesToCheck_14_7; // @[AxiLoadQueue.scala 140:26:@12207.4]
  wire  _T_13272; // @[AxiLoadQueue.scala 140:18:@12208.4]
  wire  entriesToCheck_14_8; // @[AxiLoadQueue.scala 140:26:@12209.4]
  wire  _T_13274; // @[AxiLoadQueue.scala 140:18:@12210.4]
  wire  entriesToCheck_14_9; // @[AxiLoadQueue.scala 140:26:@12211.4]
  wire  _T_13276; // @[AxiLoadQueue.scala 140:18:@12212.4]
  wire  entriesToCheck_14_10; // @[AxiLoadQueue.scala 140:26:@12213.4]
  wire  _T_13278; // @[AxiLoadQueue.scala 140:18:@12214.4]
  wire  entriesToCheck_14_11; // @[AxiLoadQueue.scala 140:26:@12215.4]
  wire  _T_13280; // @[AxiLoadQueue.scala 140:18:@12216.4]
  wire  entriesToCheck_14_12; // @[AxiLoadQueue.scala 140:26:@12217.4]
  wire  _T_13282; // @[AxiLoadQueue.scala 140:18:@12218.4]
  wire  entriesToCheck_14_13; // @[AxiLoadQueue.scala 140:26:@12219.4]
  wire  _T_13284; // @[AxiLoadQueue.scala 140:18:@12220.4]
  wire  entriesToCheck_14_14; // @[AxiLoadQueue.scala 140:26:@12221.4]
  wire  _T_13286; // @[AxiLoadQueue.scala 140:18:@12222.4]
  wire  entriesToCheck_14_15; // @[AxiLoadQueue.scala 140:26:@12223.4]
  wire  _T_13288; // @[AxiLoadQueue.scala 140:18:@12240.4]
  wire  entriesToCheck_15_0; // @[AxiLoadQueue.scala 140:26:@12241.4]
  wire  _T_13290; // @[AxiLoadQueue.scala 140:18:@12242.4]
  wire  entriesToCheck_15_1; // @[AxiLoadQueue.scala 140:26:@12243.4]
  wire  _T_13292; // @[AxiLoadQueue.scala 140:18:@12244.4]
  wire  entriesToCheck_15_2; // @[AxiLoadQueue.scala 140:26:@12245.4]
  wire  _T_13294; // @[AxiLoadQueue.scala 140:18:@12246.4]
  wire  entriesToCheck_15_3; // @[AxiLoadQueue.scala 140:26:@12247.4]
  wire  _T_13296; // @[AxiLoadQueue.scala 140:18:@12248.4]
  wire  entriesToCheck_15_4; // @[AxiLoadQueue.scala 140:26:@12249.4]
  wire  _T_13298; // @[AxiLoadQueue.scala 140:18:@12250.4]
  wire  entriesToCheck_15_5; // @[AxiLoadQueue.scala 140:26:@12251.4]
  wire  _T_13300; // @[AxiLoadQueue.scala 140:18:@12252.4]
  wire  entriesToCheck_15_6; // @[AxiLoadQueue.scala 140:26:@12253.4]
  wire  _T_13302; // @[AxiLoadQueue.scala 140:18:@12254.4]
  wire  entriesToCheck_15_7; // @[AxiLoadQueue.scala 140:26:@12255.4]
  wire  _T_13304; // @[AxiLoadQueue.scala 140:18:@12256.4]
  wire  entriesToCheck_15_8; // @[AxiLoadQueue.scala 140:26:@12257.4]
  wire  _T_13306; // @[AxiLoadQueue.scala 140:18:@12258.4]
  wire  entriesToCheck_15_9; // @[AxiLoadQueue.scala 140:26:@12259.4]
  wire  _T_13308; // @[AxiLoadQueue.scala 140:18:@12260.4]
  wire  entriesToCheck_15_10; // @[AxiLoadQueue.scala 140:26:@12261.4]
  wire  _T_13310; // @[AxiLoadQueue.scala 140:18:@12262.4]
  wire  entriesToCheck_15_11; // @[AxiLoadQueue.scala 140:26:@12263.4]
  wire  _T_13312; // @[AxiLoadQueue.scala 140:18:@12264.4]
  wire  entriesToCheck_15_12; // @[AxiLoadQueue.scala 140:26:@12265.4]
  wire  _T_13314; // @[AxiLoadQueue.scala 140:18:@12266.4]
  wire  entriesToCheck_15_13; // @[AxiLoadQueue.scala 140:26:@12267.4]
  wire  _T_13316; // @[AxiLoadQueue.scala 140:18:@12268.4]
  wire  entriesToCheck_15_14; // @[AxiLoadQueue.scala 140:26:@12269.4]
  wire  _T_13318; // @[AxiLoadQueue.scala 140:18:@12270.4]
  wire  entriesToCheck_15_15; // @[AxiLoadQueue.scala 140:26:@12271.4]
  wire  _T_14550; // @[AxiLoadQueue.scala 150:92:@12289.4]
  wire  _T_14551; // @[AxiLoadQueue.scala 151:41:@12290.4]
  wire  _T_14552; // @[AxiLoadQueue.scala 152:30:@12291.4]
  wire  conflict_0_0; // @[AxiLoadQueue.scala 151:68:@12292.4]
  wire  _T_14554; // @[AxiLoadQueue.scala 150:92:@12294.4]
  wire  _T_14555; // @[AxiLoadQueue.scala 151:41:@12295.4]
  wire  _T_14556; // @[AxiLoadQueue.scala 152:30:@12296.4]
  wire  conflict_0_1; // @[AxiLoadQueue.scala 151:68:@12297.4]
  wire  _T_14558; // @[AxiLoadQueue.scala 150:92:@12299.4]
  wire  _T_14559; // @[AxiLoadQueue.scala 151:41:@12300.4]
  wire  _T_14560; // @[AxiLoadQueue.scala 152:30:@12301.4]
  wire  conflict_0_2; // @[AxiLoadQueue.scala 151:68:@12302.4]
  wire  _T_14562; // @[AxiLoadQueue.scala 150:92:@12304.4]
  wire  _T_14563; // @[AxiLoadQueue.scala 151:41:@12305.4]
  wire  _T_14564; // @[AxiLoadQueue.scala 152:30:@12306.4]
  wire  conflict_0_3; // @[AxiLoadQueue.scala 151:68:@12307.4]
  wire  _T_14566; // @[AxiLoadQueue.scala 150:92:@12309.4]
  wire  _T_14567; // @[AxiLoadQueue.scala 151:41:@12310.4]
  wire  _T_14568; // @[AxiLoadQueue.scala 152:30:@12311.4]
  wire  conflict_0_4; // @[AxiLoadQueue.scala 151:68:@12312.4]
  wire  _T_14570; // @[AxiLoadQueue.scala 150:92:@12314.4]
  wire  _T_14571; // @[AxiLoadQueue.scala 151:41:@12315.4]
  wire  _T_14572; // @[AxiLoadQueue.scala 152:30:@12316.4]
  wire  conflict_0_5; // @[AxiLoadQueue.scala 151:68:@12317.4]
  wire  _T_14574; // @[AxiLoadQueue.scala 150:92:@12319.4]
  wire  _T_14575; // @[AxiLoadQueue.scala 151:41:@12320.4]
  wire  _T_14576; // @[AxiLoadQueue.scala 152:30:@12321.4]
  wire  conflict_0_6; // @[AxiLoadQueue.scala 151:68:@12322.4]
  wire  _T_14578; // @[AxiLoadQueue.scala 150:92:@12324.4]
  wire  _T_14579; // @[AxiLoadQueue.scala 151:41:@12325.4]
  wire  _T_14580; // @[AxiLoadQueue.scala 152:30:@12326.4]
  wire  conflict_0_7; // @[AxiLoadQueue.scala 151:68:@12327.4]
  wire  _T_14582; // @[AxiLoadQueue.scala 150:92:@12329.4]
  wire  _T_14583; // @[AxiLoadQueue.scala 151:41:@12330.4]
  wire  _T_14584; // @[AxiLoadQueue.scala 152:30:@12331.4]
  wire  conflict_0_8; // @[AxiLoadQueue.scala 151:68:@12332.4]
  wire  _T_14586; // @[AxiLoadQueue.scala 150:92:@12334.4]
  wire  _T_14587; // @[AxiLoadQueue.scala 151:41:@12335.4]
  wire  _T_14588; // @[AxiLoadQueue.scala 152:30:@12336.4]
  wire  conflict_0_9; // @[AxiLoadQueue.scala 151:68:@12337.4]
  wire  _T_14590; // @[AxiLoadQueue.scala 150:92:@12339.4]
  wire  _T_14591; // @[AxiLoadQueue.scala 151:41:@12340.4]
  wire  _T_14592; // @[AxiLoadQueue.scala 152:30:@12341.4]
  wire  conflict_0_10; // @[AxiLoadQueue.scala 151:68:@12342.4]
  wire  _T_14594; // @[AxiLoadQueue.scala 150:92:@12344.4]
  wire  _T_14595; // @[AxiLoadQueue.scala 151:41:@12345.4]
  wire  _T_14596; // @[AxiLoadQueue.scala 152:30:@12346.4]
  wire  conflict_0_11; // @[AxiLoadQueue.scala 151:68:@12347.4]
  wire  _T_14598; // @[AxiLoadQueue.scala 150:92:@12349.4]
  wire  _T_14599; // @[AxiLoadQueue.scala 151:41:@12350.4]
  wire  _T_14600; // @[AxiLoadQueue.scala 152:30:@12351.4]
  wire  conflict_0_12; // @[AxiLoadQueue.scala 151:68:@12352.4]
  wire  _T_14602; // @[AxiLoadQueue.scala 150:92:@12354.4]
  wire  _T_14603; // @[AxiLoadQueue.scala 151:41:@12355.4]
  wire  _T_14604; // @[AxiLoadQueue.scala 152:30:@12356.4]
  wire  conflict_0_13; // @[AxiLoadQueue.scala 151:68:@12357.4]
  wire  _T_14606; // @[AxiLoadQueue.scala 150:92:@12359.4]
  wire  _T_14607; // @[AxiLoadQueue.scala 151:41:@12360.4]
  wire  _T_14608; // @[AxiLoadQueue.scala 152:30:@12361.4]
  wire  conflict_0_14; // @[AxiLoadQueue.scala 151:68:@12362.4]
  wire  _T_14610; // @[AxiLoadQueue.scala 150:92:@12364.4]
  wire  _T_14611; // @[AxiLoadQueue.scala 151:41:@12365.4]
  wire  _T_14612; // @[AxiLoadQueue.scala 152:30:@12366.4]
  wire  conflict_0_15; // @[AxiLoadQueue.scala 151:68:@12367.4]
  wire  _T_14614; // @[AxiLoadQueue.scala 150:92:@12369.4]
  wire  _T_14615; // @[AxiLoadQueue.scala 151:41:@12370.4]
  wire  _T_14616; // @[AxiLoadQueue.scala 152:30:@12371.4]
  wire  conflict_1_0; // @[AxiLoadQueue.scala 151:68:@12372.4]
  wire  _T_14618; // @[AxiLoadQueue.scala 150:92:@12374.4]
  wire  _T_14619; // @[AxiLoadQueue.scala 151:41:@12375.4]
  wire  _T_14620; // @[AxiLoadQueue.scala 152:30:@12376.4]
  wire  conflict_1_1; // @[AxiLoadQueue.scala 151:68:@12377.4]
  wire  _T_14622; // @[AxiLoadQueue.scala 150:92:@12379.4]
  wire  _T_14623; // @[AxiLoadQueue.scala 151:41:@12380.4]
  wire  _T_14624; // @[AxiLoadQueue.scala 152:30:@12381.4]
  wire  conflict_1_2; // @[AxiLoadQueue.scala 151:68:@12382.4]
  wire  _T_14626; // @[AxiLoadQueue.scala 150:92:@12384.4]
  wire  _T_14627; // @[AxiLoadQueue.scala 151:41:@12385.4]
  wire  _T_14628; // @[AxiLoadQueue.scala 152:30:@12386.4]
  wire  conflict_1_3; // @[AxiLoadQueue.scala 151:68:@12387.4]
  wire  _T_14630; // @[AxiLoadQueue.scala 150:92:@12389.4]
  wire  _T_14631; // @[AxiLoadQueue.scala 151:41:@12390.4]
  wire  _T_14632; // @[AxiLoadQueue.scala 152:30:@12391.4]
  wire  conflict_1_4; // @[AxiLoadQueue.scala 151:68:@12392.4]
  wire  _T_14634; // @[AxiLoadQueue.scala 150:92:@12394.4]
  wire  _T_14635; // @[AxiLoadQueue.scala 151:41:@12395.4]
  wire  _T_14636; // @[AxiLoadQueue.scala 152:30:@12396.4]
  wire  conflict_1_5; // @[AxiLoadQueue.scala 151:68:@12397.4]
  wire  _T_14638; // @[AxiLoadQueue.scala 150:92:@12399.4]
  wire  _T_14639; // @[AxiLoadQueue.scala 151:41:@12400.4]
  wire  _T_14640; // @[AxiLoadQueue.scala 152:30:@12401.4]
  wire  conflict_1_6; // @[AxiLoadQueue.scala 151:68:@12402.4]
  wire  _T_14642; // @[AxiLoadQueue.scala 150:92:@12404.4]
  wire  _T_14643; // @[AxiLoadQueue.scala 151:41:@12405.4]
  wire  _T_14644; // @[AxiLoadQueue.scala 152:30:@12406.4]
  wire  conflict_1_7; // @[AxiLoadQueue.scala 151:68:@12407.4]
  wire  _T_14646; // @[AxiLoadQueue.scala 150:92:@12409.4]
  wire  _T_14647; // @[AxiLoadQueue.scala 151:41:@12410.4]
  wire  _T_14648; // @[AxiLoadQueue.scala 152:30:@12411.4]
  wire  conflict_1_8; // @[AxiLoadQueue.scala 151:68:@12412.4]
  wire  _T_14650; // @[AxiLoadQueue.scala 150:92:@12414.4]
  wire  _T_14651; // @[AxiLoadQueue.scala 151:41:@12415.4]
  wire  _T_14652; // @[AxiLoadQueue.scala 152:30:@12416.4]
  wire  conflict_1_9; // @[AxiLoadQueue.scala 151:68:@12417.4]
  wire  _T_14654; // @[AxiLoadQueue.scala 150:92:@12419.4]
  wire  _T_14655; // @[AxiLoadQueue.scala 151:41:@12420.4]
  wire  _T_14656; // @[AxiLoadQueue.scala 152:30:@12421.4]
  wire  conflict_1_10; // @[AxiLoadQueue.scala 151:68:@12422.4]
  wire  _T_14658; // @[AxiLoadQueue.scala 150:92:@12424.4]
  wire  _T_14659; // @[AxiLoadQueue.scala 151:41:@12425.4]
  wire  _T_14660; // @[AxiLoadQueue.scala 152:30:@12426.4]
  wire  conflict_1_11; // @[AxiLoadQueue.scala 151:68:@12427.4]
  wire  _T_14662; // @[AxiLoadQueue.scala 150:92:@12429.4]
  wire  _T_14663; // @[AxiLoadQueue.scala 151:41:@12430.4]
  wire  _T_14664; // @[AxiLoadQueue.scala 152:30:@12431.4]
  wire  conflict_1_12; // @[AxiLoadQueue.scala 151:68:@12432.4]
  wire  _T_14666; // @[AxiLoadQueue.scala 150:92:@12434.4]
  wire  _T_14667; // @[AxiLoadQueue.scala 151:41:@12435.4]
  wire  _T_14668; // @[AxiLoadQueue.scala 152:30:@12436.4]
  wire  conflict_1_13; // @[AxiLoadQueue.scala 151:68:@12437.4]
  wire  _T_14670; // @[AxiLoadQueue.scala 150:92:@12439.4]
  wire  _T_14671; // @[AxiLoadQueue.scala 151:41:@12440.4]
  wire  _T_14672; // @[AxiLoadQueue.scala 152:30:@12441.4]
  wire  conflict_1_14; // @[AxiLoadQueue.scala 151:68:@12442.4]
  wire  _T_14674; // @[AxiLoadQueue.scala 150:92:@12444.4]
  wire  _T_14675; // @[AxiLoadQueue.scala 151:41:@12445.4]
  wire  _T_14676; // @[AxiLoadQueue.scala 152:30:@12446.4]
  wire  conflict_1_15; // @[AxiLoadQueue.scala 151:68:@12447.4]
  wire  _T_14678; // @[AxiLoadQueue.scala 150:92:@12449.4]
  wire  _T_14679; // @[AxiLoadQueue.scala 151:41:@12450.4]
  wire  _T_14680; // @[AxiLoadQueue.scala 152:30:@12451.4]
  wire  conflict_2_0; // @[AxiLoadQueue.scala 151:68:@12452.4]
  wire  _T_14682; // @[AxiLoadQueue.scala 150:92:@12454.4]
  wire  _T_14683; // @[AxiLoadQueue.scala 151:41:@12455.4]
  wire  _T_14684; // @[AxiLoadQueue.scala 152:30:@12456.4]
  wire  conflict_2_1; // @[AxiLoadQueue.scala 151:68:@12457.4]
  wire  _T_14686; // @[AxiLoadQueue.scala 150:92:@12459.4]
  wire  _T_14687; // @[AxiLoadQueue.scala 151:41:@12460.4]
  wire  _T_14688; // @[AxiLoadQueue.scala 152:30:@12461.4]
  wire  conflict_2_2; // @[AxiLoadQueue.scala 151:68:@12462.4]
  wire  _T_14690; // @[AxiLoadQueue.scala 150:92:@12464.4]
  wire  _T_14691; // @[AxiLoadQueue.scala 151:41:@12465.4]
  wire  _T_14692; // @[AxiLoadQueue.scala 152:30:@12466.4]
  wire  conflict_2_3; // @[AxiLoadQueue.scala 151:68:@12467.4]
  wire  _T_14694; // @[AxiLoadQueue.scala 150:92:@12469.4]
  wire  _T_14695; // @[AxiLoadQueue.scala 151:41:@12470.4]
  wire  _T_14696; // @[AxiLoadQueue.scala 152:30:@12471.4]
  wire  conflict_2_4; // @[AxiLoadQueue.scala 151:68:@12472.4]
  wire  _T_14698; // @[AxiLoadQueue.scala 150:92:@12474.4]
  wire  _T_14699; // @[AxiLoadQueue.scala 151:41:@12475.4]
  wire  _T_14700; // @[AxiLoadQueue.scala 152:30:@12476.4]
  wire  conflict_2_5; // @[AxiLoadQueue.scala 151:68:@12477.4]
  wire  _T_14702; // @[AxiLoadQueue.scala 150:92:@12479.4]
  wire  _T_14703; // @[AxiLoadQueue.scala 151:41:@12480.4]
  wire  _T_14704; // @[AxiLoadQueue.scala 152:30:@12481.4]
  wire  conflict_2_6; // @[AxiLoadQueue.scala 151:68:@12482.4]
  wire  _T_14706; // @[AxiLoadQueue.scala 150:92:@12484.4]
  wire  _T_14707; // @[AxiLoadQueue.scala 151:41:@12485.4]
  wire  _T_14708; // @[AxiLoadQueue.scala 152:30:@12486.4]
  wire  conflict_2_7; // @[AxiLoadQueue.scala 151:68:@12487.4]
  wire  _T_14710; // @[AxiLoadQueue.scala 150:92:@12489.4]
  wire  _T_14711; // @[AxiLoadQueue.scala 151:41:@12490.4]
  wire  _T_14712; // @[AxiLoadQueue.scala 152:30:@12491.4]
  wire  conflict_2_8; // @[AxiLoadQueue.scala 151:68:@12492.4]
  wire  _T_14714; // @[AxiLoadQueue.scala 150:92:@12494.4]
  wire  _T_14715; // @[AxiLoadQueue.scala 151:41:@12495.4]
  wire  _T_14716; // @[AxiLoadQueue.scala 152:30:@12496.4]
  wire  conflict_2_9; // @[AxiLoadQueue.scala 151:68:@12497.4]
  wire  _T_14718; // @[AxiLoadQueue.scala 150:92:@12499.4]
  wire  _T_14719; // @[AxiLoadQueue.scala 151:41:@12500.4]
  wire  _T_14720; // @[AxiLoadQueue.scala 152:30:@12501.4]
  wire  conflict_2_10; // @[AxiLoadQueue.scala 151:68:@12502.4]
  wire  _T_14722; // @[AxiLoadQueue.scala 150:92:@12504.4]
  wire  _T_14723; // @[AxiLoadQueue.scala 151:41:@12505.4]
  wire  _T_14724; // @[AxiLoadQueue.scala 152:30:@12506.4]
  wire  conflict_2_11; // @[AxiLoadQueue.scala 151:68:@12507.4]
  wire  _T_14726; // @[AxiLoadQueue.scala 150:92:@12509.4]
  wire  _T_14727; // @[AxiLoadQueue.scala 151:41:@12510.4]
  wire  _T_14728; // @[AxiLoadQueue.scala 152:30:@12511.4]
  wire  conflict_2_12; // @[AxiLoadQueue.scala 151:68:@12512.4]
  wire  _T_14730; // @[AxiLoadQueue.scala 150:92:@12514.4]
  wire  _T_14731; // @[AxiLoadQueue.scala 151:41:@12515.4]
  wire  _T_14732; // @[AxiLoadQueue.scala 152:30:@12516.4]
  wire  conflict_2_13; // @[AxiLoadQueue.scala 151:68:@12517.4]
  wire  _T_14734; // @[AxiLoadQueue.scala 150:92:@12519.4]
  wire  _T_14735; // @[AxiLoadQueue.scala 151:41:@12520.4]
  wire  _T_14736; // @[AxiLoadQueue.scala 152:30:@12521.4]
  wire  conflict_2_14; // @[AxiLoadQueue.scala 151:68:@12522.4]
  wire  _T_14738; // @[AxiLoadQueue.scala 150:92:@12524.4]
  wire  _T_14739; // @[AxiLoadQueue.scala 151:41:@12525.4]
  wire  _T_14740; // @[AxiLoadQueue.scala 152:30:@12526.4]
  wire  conflict_2_15; // @[AxiLoadQueue.scala 151:68:@12527.4]
  wire  _T_14742; // @[AxiLoadQueue.scala 150:92:@12529.4]
  wire  _T_14743; // @[AxiLoadQueue.scala 151:41:@12530.4]
  wire  _T_14744; // @[AxiLoadQueue.scala 152:30:@12531.4]
  wire  conflict_3_0; // @[AxiLoadQueue.scala 151:68:@12532.4]
  wire  _T_14746; // @[AxiLoadQueue.scala 150:92:@12534.4]
  wire  _T_14747; // @[AxiLoadQueue.scala 151:41:@12535.4]
  wire  _T_14748; // @[AxiLoadQueue.scala 152:30:@12536.4]
  wire  conflict_3_1; // @[AxiLoadQueue.scala 151:68:@12537.4]
  wire  _T_14750; // @[AxiLoadQueue.scala 150:92:@12539.4]
  wire  _T_14751; // @[AxiLoadQueue.scala 151:41:@12540.4]
  wire  _T_14752; // @[AxiLoadQueue.scala 152:30:@12541.4]
  wire  conflict_3_2; // @[AxiLoadQueue.scala 151:68:@12542.4]
  wire  _T_14754; // @[AxiLoadQueue.scala 150:92:@12544.4]
  wire  _T_14755; // @[AxiLoadQueue.scala 151:41:@12545.4]
  wire  _T_14756; // @[AxiLoadQueue.scala 152:30:@12546.4]
  wire  conflict_3_3; // @[AxiLoadQueue.scala 151:68:@12547.4]
  wire  _T_14758; // @[AxiLoadQueue.scala 150:92:@12549.4]
  wire  _T_14759; // @[AxiLoadQueue.scala 151:41:@12550.4]
  wire  _T_14760; // @[AxiLoadQueue.scala 152:30:@12551.4]
  wire  conflict_3_4; // @[AxiLoadQueue.scala 151:68:@12552.4]
  wire  _T_14762; // @[AxiLoadQueue.scala 150:92:@12554.4]
  wire  _T_14763; // @[AxiLoadQueue.scala 151:41:@12555.4]
  wire  _T_14764; // @[AxiLoadQueue.scala 152:30:@12556.4]
  wire  conflict_3_5; // @[AxiLoadQueue.scala 151:68:@12557.4]
  wire  _T_14766; // @[AxiLoadQueue.scala 150:92:@12559.4]
  wire  _T_14767; // @[AxiLoadQueue.scala 151:41:@12560.4]
  wire  _T_14768; // @[AxiLoadQueue.scala 152:30:@12561.4]
  wire  conflict_3_6; // @[AxiLoadQueue.scala 151:68:@12562.4]
  wire  _T_14770; // @[AxiLoadQueue.scala 150:92:@12564.4]
  wire  _T_14771; // @[AxiLoadQueue.scala 151:41:@12565.4]
  wire  _T_14772; // @[AxiLoadQueue.scala 152:30:@12566.4]
  wire  conflict_3_7; // @[AxiLoadQueue.scala 151:68:@12567.4]
  wire  _T_14774; // @[AxiLoadQueue.scala 150:92:@12569.4]
  wire  _T_14775; // @[AxiLoadQueue.scala 151:41:@12570.4]
  wire  _T_14776; // @[AxiLoadQueue.scala 152:30:@12571.4]
  wire  conflict_3_8; // @[AxiLoadQueue.scala 151:68:@12572.4]
  wire  _T_14778; // @[AxiLoadQueue.scala 150:92:@12574.4]
  wire  _T_14779; // @[AxiLoadQueue.scala 151:41:@12575.4]
  wire  _T_14780; // @[AxiLoadQueue.scala 152:30:@12576.4]
  wire  conflict_3_9; // @[AxiLoadQueue.scala 151:68:@12577.4]
  wire  _T_14782; // @[AxiLoadQueue.scala 150:92:@12579.4]
  wire  _T_14783; // @[AxiLoadQueue.scala 151:41:@12580.4]
  wire  _T_14784; // @[AxiLoadQueue.scala 152:30:@12581.4]
  wire  conflict_3_10; // @[AxiLoadQueue.scala 151:68:@12582.4]
  wire  _T_14786; // @[AxiLoadQueue.scala 150:92:@12584.4]
  wire  _T_14787; // @[AxiLoadQueue.scala 151:41:@12585.4]
  wire  _T_14788; // @[AxiLoadQueue.scala 152:30:@12586.4]
  wire  conflict_3_11; // @[AxiLoadQueue.scala 151:68:@12587.4]
  wire  _T_14790; // @[AxiLoadQueue.scala 150:92:@12589.4]
  wire  _T_14791; // @[AxiLoadQueue.scala 151:41:@12590.4]
  wire  _T_14792; // @[AxiLoadQueue.scala 152:30:@12591.4]
  wire  conflict_3_12; // @[AxiLoadQueue.scala 151:68:@12592.4]
  wire  _T_14794; // @[AxiLoadQueue.scala 150:92:@12594.4]
  wire  _T_14795; // @[AxiLoadQueue.scala 151:41:@12595.4]
  wire  _T_14796; // @[AxiLoadQueue.scala 152:30:@12596.4]
  wire  conflict_3_13; // @[AxiLoadQueue.scala 151:68:@12597.4]
  wire  _T_14798; // @[AxiLoadQueue.scala 150:92:@12599.4]
  wire  _T_14799; // @[AxiLoadQueue.scala 151:41:@12600.4]
  wire  _T_14800; // @[AxiLoadQueue.scala 152:30:@12601.4]
  wire  conflict_3_14; // @[AxiLoadQueue.scala 151:68:@12602.4]
  wire  _T_14802; // @[AxiLoadQueue.scala 150:92:@12604.4]
  wire  _T_14803; // @[AxiLoadQueue.scala 151:41:@12605.4]
  wire  _T_14804; // @[AxiLoadQueue.scala 152:30:@12606.4]
  wire  conflict_3_15; // @[AxiLoadQueue.scala 151:68:@12607.4]
  wire  _T_14806; // @[AxiLoadQueue.scala 150:92:@12609.4]
  wire  _T_14807; // @[AxiLoadQueue.scala 151:41:@12610.4]
  wire  _T_14808; // @[AxiLoadQueue.scala 152:30:@12611.4]
  wire  conflict_4_0; // @[AxiLoadQueue.scala 151:68:@12612.4]
  wire  _T_14810; // @[AxiLoadQueue.scala 150:92:@12614.4]
  wire  _T_14811; // @[AxiLoadQueue.scala 151:41:@12615.4]
  wire  _T_14812; // @[AxiLoadQueue.scala 152:30:@12616.4]
  wire  conflict_4_1; // @[AxiLoadQueue.scala 151:68:@12617.4]
  wire  _T_14814; // @[AxiLoadQueue.scala 150:92:@12619.4]
  wire  _T_14815; // @[AxiLoadQueue.scala 151:41:@12620.4]
  wire  _T_14816; // @[AxiLoadQueue.scala 152:30:@12621.4]
  wire  conflict_4_2; // @[AxiLoadQueue.scala 151:68:@12622.4]
  wire  _T_14818; // @[AxiLoadQueue.scala 150:92:@12624.4]
  wire  _T_14819; // @[AxiLoadQueue.scala 151:41:@12625.4]
  wire  _T_14820; // @[AxiLoadQueue.scala 152:30:@12626.4]
  wire  conflict_4_3; // @[AxiLoadQueue.scala 151:68:@12627.4]
  wire  _T_14822; // @[AxiLoadQueue.scala 150:92:@12629.4]
  wire  _T_14823; // @[AxiLoadQueue.scala 151:41:@12630.4]
  wire  _T_14824; // @[AxiLoadQueue.scala 152:30:@12631.4]
  wire  conflict_4_4; // @[AxiLoadQueue.scala 151:68:@12632.4]
  wire  _T_14826; // @[AxiLoadQueue.scala 150:92:@12634.4]
  wire  _T_14827; // @[AxiLoadQueue.scala 151:41:@12635.4]
  wire  _T_14828; // @[AxiLoadQueue.scala 152:30:@12636.4]
  wire  conflict_4_5; // @[AxiLoadQueue.scala 151:68:@12637.4]
  wire  _T_14830; // @[AxiLoadQueue.scala 150:92:@12639.4]
  wire  _T_14831; // @[AxiLoadQueue.scala 151:41:@12640.4]
  wire  _T_14832; // @[AxiLoadQueue.scala 152:30:@12641.4]
  wire  conflict_4_6; // @[AxiLoadQueue.scala 151:68:@12642.4]
  wire  _T_14834; // @[AxiLoadQueue.scala 150:92:@12644.4]
  wire  _T_14835; // @[AxiLoadQueue.scala 151:41:@12645.4]
  wire  _T_14836; // @[AxiLoadQueue.scala 152:30:@12646.4]
  wire  conflict_4_7; // @[AxiLoadQueue.scala 151:68:@12647.4]
  wire  _T_14838; // @[AxiLoadQueue.scala 150:92:@12649.4]
  wire  _T_14839; // @[AxiLoadQueue.scala 151:41:@12650.4]
  wire  _T_14840; // @[AxiLoadQueue.scala 152:30:@12651.4]
  wire  conflict_4_8; // @[AxiLoadQueue.scala 151:68:@12652.4]
  wire  _T_14842; // @[AxiLoadQueue.scala 150:92:@12654.4]
  wire  _T_14843; // @[AxiLoadQueue.scala 151:41:@12655.4]
  wire  _T_14844; // @[AxiLoadQueue.scala 152:30:@12656.4]
  wire  conflict_4_9; // @[AxiLoadQueue.scala 151:68:@12657.4]
  wire  _T_14846; // @[AxiLoadQueue.scala 150:92:@12659.4]
  wire  _T_14847; // @[AxiLoadQueue.scala 151:41:@12660.4]
  wire  _T_14848; // @[AxiLoadQueue.scala 152:30:@12661.4]
  wire  conflict_4_10; // @[AxiLoadQueue.scala 151:68:@12662.4]
  wire  _T_14850; // @[AxiLoadQueue.scala 150:92:@12664.4]
  wire  _T_14851; // @[AxiLoadQueue.scala 151:41:@12665.4]
  wire  _T_14852; // @[AxiLoadQueue.scala 152:30:@12666.4]
  wire  conflict_4_11; // @[AxiLoadQueue.scala 151:68:@12667.4]
  wire  _T_14854; // @[AxiLoadQueue.scala 150:92:@12669.4]
  wire  _T_14855; // @[AxiLoadQueue.scala 151:41:@12670.4]
  wire  _T_14856; // @[AxiLoadQueue.scala 152:30:@12671.4]
  wire  conflict_4_12; // @[AxiLoadQueue.scala 151:68:@12672.4]
  wire  _T_14858; // @[AxiLoadQueue.scala 150:92:@12674.4]
  wire  _T_14859; // @[AxiLoadQueue.scala 151:41:@12675.4]
  wire  _T_14860; // @[AxiLoadQueue.scala 152:30:@12676.4]
  wire  conflict_4_13; // @[AxiLoadQueue.scala 151:68:@12677.4]
  wire  _T_14862; // @[AxiLoadQueue.scala 150:92:@12679.4]
  wire  _T_14863; // @[AxiLoadQueue.scala 151:41:@12680.4]
  wire  _T_14864; // @[AxiLoadQueue.scala 152:30:@12681.4]
  wire  conflict_4_14; // @[AxiLoadQueue.scala 151:68:@12682.4]
  wire  _T_14866; // @[AxiLoadQueue.scala 150:92:@12684.4]
  wire  _T_14867; // @[AxiLoadQueue.scala 151:41:@12685.4]
  wire  _T_14868; // @[AxiLoadQueue.scala 152:30:@12686.4]
  wire  conflict_4_15; // @[AxiLoadQueue.scala 151:68:@12687.4]
  wire  _T_14870; // @[AxiLoadQueue.scala 150:92:@12689.4]
  wire  _T_14871; // @[AxiLoadQueue.scala 151:41:@12690.4]
  wire  _T_14872; // @[AxiLoadQueue.scala 152:30:@12691.4]
  wire  conflict_5_0; // @[AxiLoadQueue.scala 151:68:@12692.4]
  wire  _T_14874; // @[AxiLoadQueue.scala 150:92:@12694.4]
  wire  _T_14875; // @[AxiLoadQueue.scala 151:41:@12695.4]
  wire  _T_14876; // @[AxiLoadQueue.scala 152:30:@12696.4]
  wire  conflict_5_1; // @[AxiLoadQueue.scala 151:68:@12697.4]
  wire  _T_14878; // @[AxiLoadQueue.scala 150:92:@12699.4]
  wire  _T_14879; // @[AxiLoadQueue.scala 151:41:@12700.4]
  wire  _T_14880; // @[AxiLoadQueue.scala 152:30:@12701.4]
  wire  conflict_5_2; // @[AxiLoadQueue.scala 151:68:@12702.4]
  wire  _T_14882; // @[AxiLoadQueue.scala 150:92:@12704.4]
  wire  _T_14883; // @[AxiLoadQueue.scala 151:41:@12705.4]
  wire  _T_14884; // @[AxiLoadQueue.scala 152:30:@12706.4]
  wire  conflict_5_3; // @[AxiLoadQueue.scala 151:68:@12707.4]
  wire  _T_14886; // @[AxiLoadQueue.scala 150:92:@12709.4]
  wire  _T_14887; // @[AxiLoadQueue.scala 151:41:@12710.4]
  wire  _T_14888; // @[AxiLoadQueue.scala 152:30:@12711.4]
  wire  conflict_5_4; // @[AxiLoadQueue.scala 151:68:@12712.4]
  wire  _T_14890; // @[AxiLoadQueue.scala 150:92:@12714.4]
  wire  _T_14891; // @[AxiLoadQueue.scala 151:41:@12715.4]
  wire  _T_14892; // @[AxiLoadQueue.scala 152:30:@12716.4]
  wire  conflict_5_5; // @[AxiLoadQueue.scala 151:68:@12717.4]
  wire  _T_14894; // @[AxiLoadQueue.scala 150:92:@12719.4]
  wire  _T_14895; // @[AxiLoadQueue.scala 151:41:@12720.4]
  wire  _T_14896; // @[AxiLoadQueue.scala 152:30:@12721.4]
  wire  conflict_5_6; // @[AxiLoadQueue.scala 151:68:@12722.4]
  wire  _T_14898; // @[AxiLoadQueue.scala 150:92:@12724.4]
  wire  _T_14899; // @[AxiLoadQueue.scala 151:41:@12725.4]
  wire  _T_14900; // @[AxiLoadQueue.scala 152:30:@12726.4]
  wire  conflict_5_7; // @[AxiLoadQueue.scala 151:68:@12727.4]
  wire  _T_14902; // @[AxiLoadQueue.scala 150:92:@12729.4]
  wire  _T_14903; // @[AxiLoadQueue.scala 151:41:@12730.4]
  wire  _T_14904; // @[AxiLoadQueue.scala 152:30:@12731.4]
  wire  conflict_5_8; // @[AxiLoadQueue.scala 151:68:@12732.4]
  wire  _T_14906; // @[AxiLoadQueue.scala 150:92:@12734.4]
  wire  _T_14907; // @[AxiLoadQueue.scala 151:41:@12735.4]
  wire  _T_14908; // @[AxiLoadQueue.scala 152:30:@12736.4]
  wire  conflict_5_9; // @[AxiLoadQueue.scala 151:68:@12737.4]
  wire  _T_14910; // @[AxiLoadQueue.scala 150:92:@12739.4]
  wire  _T_14911; // @[AxiLoadQueue.scala 151:41:@12740.4]
  wire  _T_14912; // @[AxiLoadQueue.scala 152:30:@12741.4]
  wire  conflict_5_10; // @[AxiLoadQueue.scala 151:68:@12742.4]
  wire  _T_14914; // @[AxiLoadQueue.scala 150:92:@12744.4]
  wire  _T_14915; // @[AxiLoadQueue.scala 151:41:@12745.4]
  wire  _T_14916; // @[AxiLoadQueue.scala 152:30:@12746.4]
  wire  conflict_5_11; // @[AxiLoadQueue.scala 151:68:@12747.4]
  wire  _T_14918; // @[AxiLoadQueue.scala 150:92:@12749.4]
  wire  _T_14919; // @[AxiLoadQueue.scala 151:41:@12750.4]
  wire  _T_14920; // @[AxiLoadQueue.scala 152:30:@12751.4]
  wire  conflict_5_12; // @[AxiLoadQueue.scala 151:68:@12752.4]
  wire  _T_14922; // @[AxiLoadQueue.scala 150:92:@12754.4]
  wire  _T_14923; // @[AxiLoadQueue.scala 151:41:@12755.4]
  wire  _T_14924; // @[AxiLoadQueue.scala 152:30:@12756.4]
  wire  conflict_5_13; // @[AxiLoadQueue.scala 151:68:@12757.4]
  wire  _T_14926; // @[AxiLoadQueue.scala 150:92:@12759.4]
  wire  _T_14927; // @[AxiLoadQueue.scala 151:41:@12760.4]
  wire  _T_14928; // @[AxiLoadQueue.scala 152:30:@12761.4]
  wire  conflict_5_14; // @[AxiLoadQueue.scala 151:68:@12762.4]
  wire  _T_14930; // @[AxiLoadQueue.scala 150:92:@12764.4]
  wire  _T_14931; // @[AxiLoadQueue.scala 151:41:@12765.4]
  wire  _T_14932; // @[AxiLoadQueue.scala 152:30:@12766.4]
  wire  conflict_5_15; // @[AxiLoadQueue.scala 151:68:@12767.4]
  wire  _T_14934; // @[AxiLoadQueue.scala 150:92:@12769.4]
  wire  _T_14935; // @[AxiLoadQueue.scala 151:41:@12770.4]
  wire  _T_14936; // @[AxiLoadQueue.scala 152:30:@12771.4]
  wire  conflict_6_0; // @[AxiLoadQueue.scala 151:68:@12772.4]
  wire  _T_14938; // @[AxiLoadQueue.scala 150:92:@12774.4]
  wire  _T_14939; // @[AxiLoadQueue.scala 151:41:@12775.4]
  wire  _T_14940; // @[AxiLoadQueue.scala 152:30:@12776.4]
  wire  conflict_6_1; // @[AxiLoadQueue.scala 151:68:@12777.4]
  wire  _T_14942; // @[AxiLoadQueue.scala 150:92:@12779.4]
  wire  _T_14943; // @[AxiLoadQueue.scala 151:41:@12780.4]
  wire  _T_14944; // @[AxiLoadQueue.scala 152:30:@12781.4]
  wire  conflict_6_2; // @[AxiLoadQueue.scala 151:68:@12782.4]
  wire  _T_14946; // @[AxiLoadQueue.scala 150:92:@12784.4]
  wire  _T_14947; // @[AxiLoadQueue.scala 151:41:@12785.4]
  wire  _T_14948; // @[AxiLoadQueue.scala 152:30:@12786.4]
  wire  conflict_6_3; // @[AxiLoadQueue.scala 151:68:@12787.4]
  wire  _T_14950; // @[AxiLoadQueue.scala 150:92:@12789.4]
  wire  _T_14951; // @[AxiLoadQueue.scala 151:41:@12790.4]
  wire  _T_14952; // @[AxiLoadQueue.scala 152:30:@12791.4]
  wire  conflict_6_4; // @[AxiLoadQueue.scala 151:68:@12792.4]
  wire  _T_14954; // @[AxiLoadQueue.scala 150:92:@12794.4]
  wire  _T_14955; // @[AxiLoadQueue.scala 151:41:@12795.4]
  wire  _T_14956; // @[AxiLoadQueue.scala 152:30:@12796.4]
  wire  conflict_6_5; // @[AxiLoadQueue.scala 151:68:@12797.4]
  wire  _T_14958; // @[AxiLoadQueue.scala 150:92:@12799.4]
  wire  _T_14959; // @[AxiLoadQueue.scala 151:41:@12800.4]
  wire  _T_14960; // @[AxiLoadQueue.scala 152:30:@12801.4]
  wire  conflict_6_6; // @[AxiLoadQueue.scala 151:68:@12802.4]
  wire  _T_14962; // @[AxiLoadQueue.scala 150:92:@12804.4]
  wire  _T_14963; // @[AxiLoadQueue.scala 151:41:@12805.4]
  wire  _T_14964; // @[AxiLoadQueue.scala 152:30:@12806.4]
  wire  conflict_6_7; // @[AxiLoadQueue.scala 151:68:@12807.4]
  wire  _T_14966; // @[AxiLoadQueue.scala 150:92:@12809.4]
  wire  _T_14967; // @[AxiLoadQueue.scala 151:41:@12810.4]
  wire  _T_14968; // @[AxiLoadQueue.scala 152:30:@12811.4]
  wire  conflict_6_8; // @[AxiLoadQueue.scala 151:68:@12812.4]
  wire  _T_14970; // @[AxiLoadQueue.scala 150:92:@12814.4]
  wire  _T_14971; // @[AxiLoadQueue.scala 151:41:@12815.4]
  wire  _T_14972; // @[AxiLoadQueue.scala 152:30:@12816.4]
  wire  conflict_6_9; // @[AxiLoadQueue.scala 151:68:@12817.4]
  wire  _T_14974; // @[AxiLoadQueue.scala 150:92:@12819.4]
  wire  _T_14975; // @[AxiLoadQueue.scala 151:41:@12820.4]
  wire  _T_14976; // @[AxiLoadQueue.scala 152:30:@12821.4]
  wire  conflict_6_10; // @[AxiLoadQueue.scala 151:68:@12822.4]
  wire  _T_14978; // @[AxiLoadQueue.scala 150:92:@12824.4]
  wire  _T_14979; // @[AxiLoadQueue.scala 151:41:@12825.4]
  wire  _T_14980; // @[AxiLoadQueue.scala 152:30:@12826.4]
  wire  conflict_6_11; // @[AxiLoadQueue.scala 151:68:@12827.4]
  wire  _T_14982; // @[AxiLoadQueue.scala 150:92:@12829.4]
  wire  _T_14983; // @[AxiLoadQueue.scala 151:41:@12830.4]
  wire  _T_14984; // @[AxiLoadQueue.scala 152:30:@12831.4]
  wire  conflict_6_12; // @[AxiLoadQueue.scala 151:68:@12832.4]
  wire  _T_14986; // @[AxiLoadQueue.scala 150:92:@12834.4]
  wire  _T_14987; // @[AxiLoadQueue.scala 151:41:@12835.4]
  wire  _T_14988; // @[AxiLoadQueue.scala 152:30:@12836.4]
  wire  conflict_6_13; // @[AxiLoadQueue.scala 151:68:@12837.4]
  wire  _T_14990; // @[AxiLoadQueue.scala 150:92:@12839.4]
  wire  _T_14991; // @[AxiLoadQueue.scala 151:41:@12840.4]
  wire  _T_14992; // @[AxiLoadQueue.scala 152:30:@12841.4]
  wire  conflict_6_14; // @[AxiLoadQueue.scala 151:68:@12842.4]
  wire  _T_14994; // @[AxiLoadQueue.scala 150:92:@12844.4]
  wire  _T_14995; // @[AxiLoadQueue.scala 151:41:@12845.4]
  wire  _T_14996; // @[AxiLoadQueue.scala 152:30:@12846.4]
  wire  conflict_6_15; // @[AxiLoadQueue.scala 151:68:@12847.4]
  wire  _T_14998; // @[AxiLoadQueue.scala 150:92:@12849.4]
  wire  _T_14999; // @[AxiLoadQueue.scala 151:41:@12850.4]
  wire  _T_15000; // @[AxiLoadQueue.scala 152:30:@12851.4]
  wire  conflict_7_0; // @[AxiLoadQueue.scala 151:68:@12852.4]
  wire  _T_15002; // @[AxiLoadQueue.scala 150:92:@12854.4]
  wire  _T_15003; // @[AxiLoadQueue.scala 151:41:@12855.4]
  wire  _T_15004; // @[AxiLoadQueue.scala 152:30:@12856.4]
  wire  conflict_7_1; // @[AxiLoadQueue.scala 151:68:@12857.4]
  wire  _T_15006; // @[AxiLoadQueue.scala 150:92:@12859.4]
  wire  _T_15007; // @[AxiLoadQueue.scala 151:41:@12860.4]
  wire  _T_15008; // @[AxiLoadQueue.scala 152:30:@12861.4]
  wire  conflict_7_2; // @[AxiLoadQueue.scala 151:68:@12862.4]
  wire  _T_15010; // @[AxiLoadQueue.scala 150:92:@12864.4]
  wire  _T_15011; // @[AxiLoadQueue.scala 151:41:@12865.4]
  wire  _T_15012; // @[AxiLoadQueue.scala 152:30:@12866.4]
  wire  conflict_7_3; // @[AxiLoadQueue.scala 151:68:@12867.4]
  wire  _T_15014; // @[AxiLoadQueue.scala 150:92:@12869.4]
  wire  _T_15015; // @[AxiLoadQueue.scala 151:41:@12870.4]
  wire  _T_15016; // @[AxiLoadQueue.scala 152:30:@12871.4]
  wire  conflict_7_4; // @[AxiLoadQueue.scala 151:68:@12872.4]
  wire  _T_15018; // @[AxiLoadQueue.scala 150:92:@12874.4]
  wire  _T_15019; // @[AxiLoadQueue.scala 151:41:@12875.4]
  wire  _T_15020; // @[AxiLoadQueue.scala 152:30:@12876.4]
  wire  conflict_7_5; // @[AxiLoadQueue.scala 151:68:@12877.4]
  wire  _T_15022; // @[AxiLoadQueue.scala 150:92:@12879.4]
  wire  _T_15023; // @[AxiLoadQueue.scala 151:41:@12880.4]
  wire  _T_15024; // @[AxiLoadQueue.scala 152:30:@12881.4]
  wire  conflict_7_6; // @[AxiLoadQueue.scala 151:68:@12882.4]
  wire  _T_15026; // @[AxiLoadQueue.scala 150:92:@12884.4]
  wire  _T_15027; // @[AxiLoadQueue.scala 151:41:@12885.4]
  wire  _T_15028; // @[AxiLoadQueue.scala 152:30:@12886.4]
  wire  conflict_7_7; // @[AxiLoadQueue.scala 151:68:@12887.4]
  wire  _T_15030; // @[AxiLoadQueue.scala 150:92:@12889.4]
  wire  _T_15031; // @[AxiLoadQueue.scala 151:41:@12890.4]
  wire  _T_15032; // @[AxiLoadQueue.scala 152:30:@12891.4]
  wire  conflict_7_8; // @[AxiLoadQueue.scala 151:68:@12892.4]
  wire  _T_15034; // @[AxiLoadQueue.scala 150:92:@12894.4]
  wire  _T_15035; // @[AxiLoadQueue.scala 151:41:@12895.4]
  wire  _T_15036; // @[AxiLoadQueue.scala 152:30:@12896.4]
  wire  conflict_7_9; // @[AxiLoadQueue.scala 151:68:@12897.4]
  wire  _T_15038; // @[AxiLoadQueue.scala 150:92:@12899.4]
  wire  _T_15039; // @[AxiLoadQueue.scala 151:41:@12900.4]
  wire  _T_15040; // @[AxiLoadQueue.scala 152:30:@12901.4]
  wire  conflict_7_10; // @[AxiLoadQueue.scala 151:68:@12902.4]
  wire  _T_15042; // @[AxiLoadQueue.scala 150:92:@12904.4]
  wire  _T_15043; // @[AxiLoadQueue.scala 151:41:@12905.4]
  wire  _T_15044; // @[AxiLoadQueue.scala 152:30:@12906.4]
  wire  conflict_7_11; // @[AxiLoadQueue.scala 151:68:@12907.4]
  wire  _T_15046; // @[AxiLoadQueue.scala 150:92:@12909.4]
  wire  _T_15047; // @[AxiLoadQueue.scala 151:41:@12910.4]
  wire  _T_15048; // @[AxiLoadQueue.scala 152:30:@12911.4]
  wire  conflict_7_12; // @[AxiLoadQueue.scala 151:68:@12912.4]
  wire  _T_15050; // @[AxiLoadQueue.scala 150:92:@12914.4]
  wire  _T_15051; // @[AxiLoadQueue.scala 151:41:@12915.4]
  wire  _T_15052; // @[AxiLoadQueue.scala 152:30:@12916.4]
  wire  conflict_7_13; // @[AxiLoadQueue.scala 151:68:@12917.4]
  wire  _T_15054; // @[AxiLoadQueue.scala 150:92:@12919.4]
  wire  _T_15055; // @[AxiLoadQueue.scala 151:41:@12920.4]
  wire  _T_15056; // @[AxiLoadQueue.scala 152:30:@12921.4]
  wire  conflict_7_14; // @[AxiLoadQueue.scala 151:68:@12922.4]
  wire  _T_15058; // @[AxiLoadQueue.scala 150:92:@12924.4]
  wire  _T_15059; // @[AxiLoadQueue.scala 151:41:@12925.4]
  wire  _T_15060; // @[AxiLoadQueue.scala 152:30:@12926.4]
  wire  conflict_7_15; // @[AxiLoadQueue.scala 151:68:@12927.4]
  wire  _T_15062; // @[AxiLoadQueue.scala 150:92:@12929.4]
  wire  _T_15063; // @[AxiLoadQueue.scala 151:41:@12930.4]
  wire  _T_15064; // @[AxiLoadQueue.scala 152:30:@12931.4]
  wire  conflict_8_0; // @[AxiLoadQueue.scala 151:68:@12932.4]
  wire  _T_15066; // @[AxiLoadQueue.scala 150:92:@12934.4]
  wire  _T_15067; // @[AxiLoadQueue.scala 151:41:@12935.4]
  wire  _T_15068; // @[AxiLoadQueue.scala 152:30:@12936.4]
  wire  conflict_8_1; // @[AxiLoadQueue.scala 151:68:@12937.4]
  wire  _T_15070; // @[AxiLoadQueue.scala 150:92:@12939.4]
  wire  _T_15071; // @[AxiLoadQueue.scala 151:41:@12940.4]
  wire  _T_15072; // @[AxiLoadQueue.scala 152:30:@12941.4]
  wire  conflict_8_2; // @[AxiLoadQueue.scala 151:68:@12942.4]
  wire  _T_15074; // @[AxiLoadQueue.scala 150:92:@12944.4]
  wire  _T_15075; // @[AxiLoadQueue.scala 151:41:@12945.4]
  wire  _T_15076; // @[AxiLoadQueue.scala 152:30:@12946.4]
  wire  conflict_8_3; // @[AxiLoadQueue.scala 151:68:@12947.4]
  wire  _T_15078; // @[AxiLoadQueue.scala 150:92:@12949.4]
  wire  _T_15079; // @[AxiLoadQueue.scala 151:41:@12950.4]
  wire  _T_15080; // @[AxiLoadQueue.scala 152:30:@12951.4]
  wire  conflict_8_4; // @[AxiLoadQueue.scala 151:68:@12952.4]
  wire  _T_15082; // @[AxiLoadQueue.scala 150:92:@12954.4]
  wire  _T_15083; // @[AxiLoadQueue.scala 151:41:@12955.4]
  wire  _T_15084; // @[AxiLoadQueue.scala 152:30:@12956.4]
  wire  conflict_8_5; // @[AxiLoadQueue.scala 151:68:@12957.4]
  wire  _T_15086; // @[AxiLoadQueue.scala 150:92:@12959.4]
  wire  _T_15087; // @[AxiLoadQueue.scala 151:41:@12960.4]
  wire  _T_15088; // @[AxiLoadQueue.scala 152:30:@12961.4]
  wire  conflict_8_6; // @[AxiLoadQueue.scala 151:68:@12962.4]
  wire  _T_15090; // @[AxiLoadQueue.scala 150:92:@12964.4]
  wire  _T_15091; // @[AxiLoadQueue.scala 151:41:@12965.4]
  wire  _T_15092; // @[AxiLoadQueue.scala 152:30:@12966.4]
  wire  conflict_8_7; // @[AxiLoadQueue.scala 151:68:@12967.4]
  wire  _T_15094; // @[AxiLoadQueue.scala 150:92:@12969.4]
  wire  _T_15095; // @[AxiLoadQueue.scala 151:41:@12970.4]
  wire  _T_15096; // @[AxiLoadQueue.scala 152:30:@12971.4]
  wire  conflict_8_8; // @[AxiLoadQueue.scala 151:68:@12972.4]
  wire  _T_15098; // @[AxiLoadQueue.scala 150:92:@12974.4]
  wire  _T_15099; // @[AxiLoadQueue.scala 151:41:@12975.4]
  wire  _T_15100; // @[AxiLoadQueue.scala 152:30:@12976.4]
  wire  conflict_8_9; // @[AxiLoadQueue.scala 151:68:@12977.4]
  wire  _T_15102; // @[AxiLoadQueue.scala 150:92:@12979.4]
  wire  _T_15103; // @[AxiLoadQueue.scala 151:41:@12980.4]
  wire  _T_15104; // @[AxiLoadQueue.scala 152:30:@12981.4]
  wire  conflict_8_10; // @[AxiLoadQueue.scala 151:68:@12982.4]
  wire  _T_15106; // @[AxiLoadQueue.scala 150:92:@12984.4]
  wire  _T_15107; // @[AxiLoadQueue.scala 151:41:@12985.4]
  wire  _T_15108; // @[AxiLoadQueue.scala 152:30:@12986.4]
  wire  conflict_8_11; // @[AxiLoadQueue.scala 151:68:@12987.4]
  wire  _T_15110; // @[AxiLoadQueue.scala 150:92:@12989.4]
  wire  _T_15111; // @[AxiLoadQueue.scala 151:41:@12990.4]
  wire  _T_15112; // @[AxiLoadQueue.scala 152:30:@12991.4]
  wire  conflict_8_12; // @[AxiLoadQueue.scala 151:68:@12992.4]
  wire  _T_15114; // @[AxiLoadQueue.scala 150:92:@12994.4]
  wire  _T_15115; // @[AxiLoadQueue.scala 151:41:@12995.4]
  wire  _T_15116; // @[AxiLoadQueue.scala 152:30:@12996.4]
  wire  conflict_8_13; // @[AxiLoadQueue.scala 151:68:@12997.4]
  wire  _T_15118; // @[AxiLoadQueue.scala 150:92:@12999.4]
  wire  _T_15119; // @[AxiLoadQueue.scala 151:41:@13000.4]
  wire  _T_15120; // @[AxiLoadQueue.scala 152:30:@13001.4]
  wire  conflict_8_14; // @[AxiLoadQueue.scala 151:68:@13002.4]
  wire  _T_15122; // @[AxiLoadQueue.scala 150:92:@13004.4]
  wire  _T_15123; // @[AxiLoadQueue.scala 151:41:@13005.4]
  wire  _T_15124; // @[AxiLoadQueue.scala 152:30:@13006.4]
  wire  conflict_8_15; // @[AxiLoadQueue.scala 151:68:@13007.4]
  wire  _T_15126; // @[AxiLoadQueue.scala 150:92:@13009.4]
  wire  _T_15127; // @[AxiLoadQueue.scala 151:41:@13010.4]
  wire  _T_15128; // @[AxiLoadQueue.scala 152:30:@13011.4]
  wire  conflict_9_0; // @[AxiLoadQueue.scala 151:68:@13012.4]
  wire  _T_15130; // @[AxiLoadQueue.scala 150:92:@13014.4]
  wire  _T_15131; // @[AxiLoadQueue.scala 151:41:@13015.4]
  wire  _T_15132; // @[AxiLoadQueue.scala 152:30:@13016.4]
  wire  conflict_9_1; // @[AxiLoadQueue.scala 151:68:@13017.4]
  wire  _T_15134; // @[AxiLoadQueue.scala 150:92:@13019.4]
  wire  _T_15135; // @[AxiLoadQueue.scala 151:41:@13020.4]
  wire  _T_15136; // @[AxiLoadQueue.scala 152:30:@13021.4]
  wire  conflict_9_2; // @[AxiLoadQueue.scala 151:68:@13022.4]
  wire  _T_15138; // @[AxiLoadQueue.scala 150:92:@13024.4]
  wire  _T_15139; // @[AxiLoadQueue.scala 151:41:@13025.4]
  wire  _T_15140; // @[AxiLoadQueue.scala 152:30:@13026.4]
  wire  conflict_9_3; // @[AxiLoadQueue.scala 151:68:@13027.4]
  wire  _T_15142; // @[AxiLoadQueue.scala 150:92:@13029.4]
  wire  _T_15143; // @[AxiLoadQueue.scala 151:41:@13030.4]
  wire  _T_15144; // @[AxiLoadQueue.scala 152:30:@13031.4]
  wire  conflict_9_4; // @[AxiLoadQueue.scala 151:68:@13032.4]
  wire  _T_15146; // @[AxiLoadQueue.scala 150:92:@13034.4]
  wire  _T_15147; // @[AxiLoadQueue.scala 151:41:@13035.4]
  wire  _T_15148; // @[AxiLoadQueue.scala 152:30:@13036.4]
  wire  conflict_9_5; // @[AxiLoadQueue.scala 151:68:@13037.4]
  wire  _T_15150; // @[AxiLoadQueue.scala 150:92:@13039.4]
  wire  _T_15151; // @[AxiLoadQueue.scala 151:41:@13040.4]
  wire  _T_15152; // @[AxiLoadQueue.scala 152:30:@13041.4]
  wire  conflict_9_6; // @[AxiLoadQueue.scala 151:68:@13042.4]
  wire  _T_15154; // @[AxiLoadQueue.scala 150:92:@13044.4]
  wire  _T_15155; // @[AxiLoadQueue.scala 151:41:@13045.4]
  wire  _T_15156; // @[AxiLoadQueue.scala 152:30:@13046.4]
  wire  conflict_9_7; // @[AxiLoadQueue.scala 151:68:@13047.4]
  wire  _T_15158; // @[AxiLoadQueue.scala 150:92:@13049.4]
  wire  _T_15159; // @[AxiLoadQueue.scala 151:41:@13050.4]
  wire  _T_15160; // @[AxiLoadQueue.scala 152:30:@13051.4]
  wire  conflict_9_8; // @[AxiLoadQueue.scala 151:68:@13052.4]
  wire  _T_15162; // @[AxiLoadQueue.scala 150:92:@13054.4]
  wire  _T_15163; // @[AxiLoadQueue.scala 151:41:@13055.4]
  wire  _T_15164; // @[AxiLoadQueue.scala 152:30:@13056.4]
  wire  conflict_9_9; // @[AxiLoadQueue.scala 151:68:@13057.4]
  wire  _T_15166; // @[AxiLoadQueue.scala 150:92:@13059.4]
  wire  _T_15167; // @[AxiLoadQueue.scala 151:41:@13060.4]
  wire  _T_15168; // @[AxiLoadQueue.scala 152:30:@13061.4]
  wire  conflict_9_10; // @[AxiLoadQueue.scala 151:68:@13062.4]
  wire  _T_15170; // @[AxiLoadQueue.scala 150:92:@13064.4]
  wire  _T_15171; // @[AxiLoadQueue.scala 151:41:@13065.4]
  wire  _T_15172; // @[AxiLoadQueue.scala 152:30:@13066.4]
  wire  conflict_9_11; // @[AxiLoadQueue.scala 151:68:@13067.4]
  wire  _T_15174; // @[AxiLoadQueue.scala 150:92:@13069.4]
  wire  _T_15175; // @[AxiLoadQueue.scala 151:41:@13070.4]
  wire  _T_15176; // @[AxiLoadQueue.scala 152:30:@13071.4]
  wire  conflict_9_12; // @[AxiLoadQueue.scala 151:68:@13072.4]
  wire  _T_15178; // @[AxiLoadQueue.scala 150:92:@13074.4]
  wire  _T_15179; // @[AxiLoadQueue.scala 151:41:@13075.4]
  wire  _T_15180; // @[AxiLoadQueue.scala 152:30:@13076.4]
  wire  conflict_9_13; // @[AxiLoadQueue.scala 151:68:@13077.4]
  wire  _T_15182; // @[AxiLoadQueue.scala 150:92:@13079.4]
  wire  _T_15183; // @[AxiLoadQueue.scala 151:41:@13080.4]
  wire  _T_15184; // @[AxiLoadQueue.scala 152:30:@13081.4]
  wire  conflict_9_14; // @[AxiLoadQueue.scala 151:68:@13082.4]
  wire  _T_15186; // @[AxiLoadQueue.scala 150:92:@13084.4]
  wire  _T_15187; // @[AxiLoadQueue.scala 151:41:@13085.4]
  wire  _T_15188; // @[AxiLoadQueue.scala 152:30:@13086.4]
  wire  conflict_9_15; // @[AxiLoadQueue.scala 151:68:@13087.4]
  wire  _T_15190; // @[AxiLoadQueue.scala 150:92:@13089.4]
  wire  _T_15191; // @[AxiLoadQueue.scala 151:41:@13090.4]
  wire  _T_15192; // @[AxiLoadQueue.scala 152:30:@13091.4]
  wire  conflict_10_0; // @[AxiLoadQueue.scala 151:68:@13092.4]
  wire  _T_15194; // @[AxiLoadQueue.scala 150:92:@13094.4]
  wire  _T_15195; // @[AxiLoadQueue.scala 151:41:@13095.4]
  wire  _T_15196; // @[AxiLoadQueue.scala 152:30:@13096.4]
  wire  conflict_10_1; // @[AxiLoadQueue.scala 151:68:@13097.4]
  wire  _T_15198; // @[AxiLoadQueue.scala 150:92:@13099.4]
  wire  _T_15199; // @[AxiLoadQueue.scala 151:41:@13100.4]
  wire  _T_15200; // @[AxiLoadQueue.scala 152:30:@13101.4]
  wire  conflict_10_2; // @[AxiLoadQueue.scala 151:68:@13102.4]
  wire  _T_15202; // @[AxiLoadQueue.scala 150:92:@13104.4]
  wire  _T_15203; // @[AxiLoadQueue.scala 151:41:@13105.4]
  wire  _T_15204; // @[AxiLoadQueue.scala 152:30:@13106.4]
  wire  conflict_10_3; // @[AxiLoadQueue.scala 151:68:@13107.4]
  wire  _T_15206; // @[AxiLoadQueue.scala 150:92:@13109.4]
  wire  _T_15207; // @[AxiLoadQueue.scala 151:41:@13110.4]
  wire  _T_15208; // @[AxiLoadQueue.scala 152:30:@13111.4]
  wire  conflict_10_4; // @[AxiLoadQueue.scala 151:68:@13112.4]
  wire  _T_15210; // @[AxiLoadQueue.scala 150:92:@13114.4]
  wire  _T_15211; // @[AxiLoadQueue.scala 151:41:@13115.4]
  wire  _T_15212; // @[AxiLoadQueue.scala 152:30:@13116.4]
  wire  conflict_10_5; // @[AxiLoadQueue.scala 151:68:@13117.4]
  wire  _T_15214; // @[AxiLoadQueue.scala 150:92:@13119.4]
  wire  _T_15215; // @[AxiLoadQueue.scala 151:41:@13120.4]
  wire  _T_15216; // @[AxiLoadQueue.scala 152:30:@13121.4]
  wire  conflict_10_6; // @[AxiLoadQueue.scala 151:68:@13122.4]
  wire  _T_15218; // @[AxiLoadQueue.scala 150:92:@13124.4]
  wire  _T_15219; // @[AxiLoadQueue.scala 151:41:@13125.4]
  wire  _T_15220; // @[AxiLoadQueue.scala 152:30:@13126.4]
  wire  conflict_10_7; // @[AxiLoadQueue.scala 151:68:@13127.4]
  wire  _T_15222; // @[AxiLoadQueue.scala 150:92:@13129.4]
  wire  _T_15223; // @[AxiLoadQueue.scala 151:41:@13130.4]
  wire  _T_15224; // @[AxiLoadQueue.scala 152:30:@13131.4]
  wire  conflict_10_8; // @[AxiLoadQueue.scala 151:68:@13132.4]
  wire  _T_15226; // @[AxiLoadQueue.scala 150:92:@13134.4]
  wire  _T_15227; // @[AxiLoadQueue.scala 151:41:@13135.4]
  wire  _T_15228; // @[AxiLoadQueue.scala 152:30:@13136.4]
  wire  conflict_10_9; // @[AxiLoadQueue.scala 151:68:@13137.4]
  wire  _T_15230; // @[AxiLoadQueue.scala 150:92:@13139.4]
  wire  _T_15231; // @[AxiLoadQueue.scala 151:41:@13140.4]
  wire  _T_15232; // @[AxiLoadQueue.scala 152:30:@13141.4]
  wire  conflict_10_10; // @[AxiLoadQueue.scala 151:68:@13142.4]
  wire  _T_15234; // @[AxiLoadQueue.scala 150:92:@13144.4]
  wire  _T_15235; // @[AxiLoadQueue.scala 151:41:@13145.4]
  wire  _T_15236; // @[AxiLoadQueue.scala 152:30:@13146.4]
  wire  conflict_10_11; // @[AxiLoadQueue.scala 151:68:@13147.4]
  wire  _T_15238; // @[AxiLoadQueue.scala 150:92:@13149.4]
  wire  _T_15239; // @[AxiLoadQueue.scala 151:41:@13150.4]
  wire  _T_15240; // @[AxiLoadQueue.scala 152:30:@13151.4]
  wire  conflict_10_12; // @[AxiLoadQueue.scala 151:68:@13152.4]
  wire  _T_15242; // @[AxiLoadQueue.scala 150:92:@13154.4]
  wire  _T_15243; // @[AxiLoadQueue.scala 151:41:@13155.4]
  wire  _T_15244; // @[AxiLoadQueue.scala 152:30:@13156.4]
  wire  conflict_10_13; // @[AxiLoadQueue.scala 151:68:@13157.4]
  wire  _T_15246; // @[AxiLoadQueue.scala 150:92:@13159.4]
  wire  _T_15247; // @[AxiLoadQueue.scala 151:41:@13160.4]
  wire  _T_15248; // @[AxiLoadQueue.scala 152:30:@13161.4]
  wire  conflict_10_14; // @[AxiLoadQueue.scala 151:68:@13162.4]
  wire  _T_15250; // @[AxiLoadQueue.scala 150:92:@13164.4]
  wire  _T_15251; // @[AxiLoadQueue.scala 151:41:@13165.4]
  wire  _T_15252; // @[AxiLoadQueue.scala 152:30:@13166.4]
  wire  conflict_10_15; // @[AxiLoadQueue.scala 151:68:@13167.4]
  wire  _T_15254; // @[AxiLoadQueue.scala 150:92:@13169.4]
  wire  _T_15255; // @[AxiLoadQueue.scala 151:41:@13170.4]
  wire  _T_15256; // @[AxiLoadQueue.scala 152:30:@13171.4]
  wire  conflict_11_0; // @[AxiLoadQueue.scala 151:68:@13172.4]
  wire  _T_15258; // @[AxiLoadQueue.scala 150:92:@13174.4]
  wire  _T_15259; // @[AxiLoadQueue.scala 151:41:@13175.4]
  wire  _T_15260; // @[AxiLoadQueue.scala 152:30:@13176.4]
  wire  conflict_11_1; // @[AxiLoadQueue.scala 151:68:@13177.4]
  wire  _T_15262; // @[AxiLoadQueue.scala 150:92:@13179.4]
  wire  _T_15263; // @[AxiLoadQueue.scala 151:41:@13180.4]
  wire  _T_15264; // @[AxiLoadQueue.scala 152:30:@13181.4]
  wire  conflict_11_2; // @[AxiLoadQueue.scala 151:68:@13182.4]
  wire  _T_15266; // @[AxiLoadQueue.scala 150:92:@13184.4]
  wire  _T_15267; // @[AxiLoadQueue.scala 151:41:@13185.4]
  wire  _T_15268; // @[AxiLoadQueue.scala 152:30:@13186.4]
  wire  conflict_11_3; // @[AxiLoadQueue.scala 151:68:@13187.4]
  wire  _T_15270; // @[AxiLoadQueue.scala 150:92:@13189.4]
  wire  _T_15271; // @[AxiLoadQueue.scala 151:41:@13190.4]
  wire  _T_15272; // @[AxiLoadQueue.scala 152:30:@13191.4]
  wire  conflict_11_4; // @[AxiLoadQueue.scala 151:68:@13192.4]
  wire  _T_15274; // @[AxiLoadQueue.scala 150:92:@13194.4]
  wire  _T_15275; // @[AxiLoadQueue.scala 151:41:@13195.4]
  wire  _T_15276; // @[AxiLoadQueue.scala 152:30:@13196.4]
  wire  conflict_11_5; // @[AxiLoadQueue.scala 151:68:@13197.4]
  wire  _T_15278; // @[AxiLoadQueue.scala 150:92:@13199.4]
  wire  _T_15279; // @[AxiLoadQueue.scala 151:41:@13200.4]
  wire  _T_15280; // @[AxiLoadQueue.scala 152:30:@13201.4]
  wire  conflict_11_6; // @[AxiLoadQueue.scala 151:68:@13202.4]
  wire  _T_15282; // @[AxiLoadQueue.scala 150:92:@13204.4]
  wire  _T_15283; // @[AxiLoadQueue.scala 151:41:@13205.4]
  wire  _T_15284; // @[AxiLoadQueue.scala 152:30:@13206.4]
  wire  conflict_11_7; // @[AxiLoadQueue.scala 151:68:@13207.4]
  wire  _T_15286; // @[AxiLoadQueue.scala 150:92:@13209.4]
  wire  _T_15287; // @[AxiLoadQueue.scala 151:41:@13210.4]
  wire  _T_15288; // @[AxiLoadQueue.scala 152:30:@13211.4]
  wire  conflict_11_8; // @[AxiLoadQueue.scala 151:68:@13212.4]
  wire  _T_15290; // @[AxiLoadQueue.scala 150:92:@13214.4]
  wire  _T_15291; // @[AxiLoadQueue.scala 151:41:@13215.4]
  wire  _T_15292; // @[AxiLoadQueue.scala 152:30:@13216.4]
  wire  conflict_11_9; // @[AxiLoadQueue.scala 151:68:@13217.4]
  wire  _T_15294; // @[AxiLoadQueue.scala 150:92:@13219.4]
  wire  _T_15295; // @[AxiLoadQueue.scala 151:41:@13220.4]
  wire  _T_15296; // @[AxiLoadQueue.scala 152:30:@13221.4]
  wire  conflict_11_10; // @[AxiLoadQueue.scala 151:68:@13222.4]
  wire  _T_15298; // @[AxiLoadQueue.scala 150:92:@13224.4]
  wire  _T_15299; // @[AxiLoadQueue.scala 151:41:@13225.4]
  wire  _T_15300; // @[AxiLoadQueue.scala 152:30:@13226.4]
  wire  conflict_11_11; // @[AxiLoadQueue.scala 151:68:@13227.4]
  wire  _T_15302; // @[AxiLoadQueue.scala 150:92:@13229.4]
  wire  _T_15303; // @[AxiLoadQueue.scala 151:41:@13230.4]
  wire  _T_15304; // @[AxiLoadQueue.scala 152:30:@13231.4]
  wire  conflict_11_12; // @[AxiLoadQueue.scala 151:68:@13232.4]
  wire  _T_15306; // @[AxiLoadQueue.scala 150:92:@13234.4]
  wire  _T_15307; // @[AxiLoadQueue.scala 151:41:@13235.4]
  wire  _T_15308; // @[AxiLoadQueue.scala 152:30:@13236.4]
  wire  conflict_11_13; // @[AxiLoadQueue.scala 151:68:@13237.4]
  wire  _T_15310; // @[AxiLoadQueue.scala 150:92:@13239.4]
  wire  _T_15311; // @[AxiLoadQueue.scala 151:41:@13240.4]
  wire  _T_15312; // @[AxiLoadQueue.scala 152:30:@13241.4]
  wire  conflict_11_14; // @[AxiLoadQueue.scala 151:68:@13242.4]
  wire  _T_15314; // @[AxiLoadQueue.scala 150:92:@13244.4]
  wire  _T_15315; // @[AxiLoadQueue.scala 151:41:@13245.4]
  wire  _T_15316; // @[AxiLoadQueue.scala 152:30:@13246.4]
  wire  conflict_11_15; // @[AxiLoadQueue.scala 151:68:@13247.4]
  wire  _T_15318; // @[AxiLoadQueue.scala 150:92:@13249.4]
  wire  _T_15319; // @[AxiLoadQueue.scala 151:41:@13250.4]
  wire  _T_15320; // @[AxiLoadQueue.scala 152:30:@13251.4]
  wire  conflict_12_0; // @[AxiLoadQueue.scala 151:68:@13252.4]
  wire  _T_15322; // @[AxiLoadQueue.scala 150:92:@13254.4]
  wire  _T_15323; // @[AxiLoadQueue.scala 151:41:@13255.4]
  wire  _T_15324; // @[AxiLoadQueue.scala 152:30:@13256.4]
  wire  conflict_12_1; // @[AxiLoadQueue.scala 151:68:@13257.4]
  wire  _T_15326; // @[AxiLoadQueue.scala 150:92:@13259.4]
  wire  _T_15327; // @[AxiLoadQueue.scala 151:41:@13260.4]
  wire  _T_15328; // @[AxiLoadQueue.scala 152:30:@13261.4]
  wire  conflict_12_2; // @[AxiLoadQueue.scala 151:68:@13262.4]
  wire  _T_15330; // @[AxiLoadQueue.scala 150:92:@13264.4]
  wire  _T_15331; // @[AxiLoadQueue.scala 151:41:@13265.4]
  wire  _T_15332; // @[AxiLoadQueue.scala 152:30:@13266.4]
  wire  conflict_12_3; // @[AxiLoadQueue.scala 151:68:@13267.4]
  wire  _T_15334; // @[AxiLoadQueue.scala 150:92:@13269.4]
  wire  _T_15335; // @[AxiLoadQueue.scala 151:41:@13270.4]
  wire  _T_15336; // @[AxiLoadQueue.scala 152:30:@13271.4]
  wire  conflict_12_4; // @[AxiLoadQueue.scala 151:68:@13272.4]
  wire  _T_15338; // @[AxiLoadQueue.scala 150:92:@13274.4]
  wire  _T_15339; // @[AxiLoadQueue.scala 151:41:@13275.4]
  wire  _T_15340; // @[AxiLoadQueue.scala 152:30:@13276.4]
  wire  conflict_12_5; // @[AxiLoadQueue.scala 151:68:@13277.4]
  wire  _T_15342; // @[AxiLoadQueue.scala 150:92:@13279.4]
  wire  _T_15343; // @[AxiLoadQueue.scala 151:41:@13280.4]
  wire  _T_15344; // @[AxiLoadQueue.scala 152:30:@13281.4]
  wire  conflict_12_6; // @[AxiLoadQueue.scala 151:68:@13282.4]
  wire  _T_15346; // @[AxiLoadQueue.scala 150:92:@13284.4]
  wire  _T_15347; // @[AxiLoadQueue.scala 151:41:@13285.4]
  wire  _T_15348; // @[AxiLoadQueue.scala 152:30:@13286.4]
  wire  conflict_12_7; // @[AxiLoadQueue.scala 151:68:@13287.4]
  wire  _T_15350; // @[AxiLoadQueue.scala 150:92:@13289.4]
  wire  _T_15351; // @[AxiLoadQueue.scala 151:41:@13290.4]
  wire  _T_15352; // @[AxiLoadQueue.scala 152:30:@13291.4]
  wire  conflict_12_8; // @[AxiLoadQueue.scala 151:68:@13292.4]
  wire  _T_15354; // @[AxiLoadQueue.scala 150:92:@13294.4]
  wire  _T_15355; // @[AxiLoadQueue.scala 151:41:@13295.4]
  wire  _T_15356; // @[AxiLoadQueue.scala 152:30:@13296.4]
  wire  conflict_12_9; // @[AxiLoadQueue.scala 151:68:@13297.4]
  wire  _T_15358; // @[AxiLoadQueue.scala 150:92:@13299.4]
  wire  _T_15359; // @[AxiLoadQueue.scala 151:41:@13300.4]
  wire  _T_15360; // @[AxiLoadQueue.scala 152:30:@13301.4]
  wire  conflict_12_10; // @[AxiLoadQueue.scala 151:68:@13302.4]
  wire  _T_15362; // @[AxiLoadQueue.scala 150:92:@13304.4]
  wire  _T_15363; // @[AxiLoadQueue.scala 151:41:@13305.4]
  wire  _T_15364; // @[AxiLoadQueue.scala 152:30:@13306.4]
  wire  conflict_12_11; // @[AxiLoadQueue.scala 151:68:@13307.4]
  wire  _T_15366; // @[AxiLoadQueue.scala 150:92:@13309.4]
  wire  _T_15367; // @[AxiLoadQueue.scala 151:41:@13310.4]
  wire  _T_15368; // @[AxiLoadQueue.scala 152:30:@13311.4]
  wire  conflict_12_12; // @[AxiLoadQueue.scala 151:68:@13312.4]
  wire  _T_15370; // @[AxiLoadQueue.scala 150:92:@13314.4]
  wire  _T_15371; // @[AxiLoadQueue.scala 151:41:@13315.4]
  wire  _T_15372; // @[AxiLoadQueue.scala 152:30:@13316.4]
  wire  conflict_12_13; // @[AxiLoadQueue.scala 151:68:@13317.4]
  wire  _T_15374; // @[AxiLoadQueue.scala 150:92:@13319.4]
  wire  _T_15375; // @[AxiLoadQueue.scala 151:41:@13320.4]
  wire  _T_15376; // @[AxiLoadQueue.scala 152:30:@13321.4]
  wire  conflict_12_14; // @[AxiLoadQueue.scala 151:68:@13322.4]
  wire  _T_15378; // @[AxiLoadQueue.scala 150:92:@13324.4]
  wire  _T_15379; // @[AxiLoadQueue.scala 151:41:@13325.4]
  wire  _T_15380; // @[AxiLoadQueue.scala 152:30:@13326.4]
  wire  conflict_12_15; // @[AxiLoadQueue.scala 151:68:@13327.4]
  wire  _T_15382; // @[AxiLoadQueue.scala 150:92:@13329.4]
  wire  _T_15383; // @[AxiLoadQueue.scala 151:41:@13330.4]
  wire  _T_15384; // @[AxiLoadQueue.scala 152:30:@13331.4]
  wire  conflict_13_0; // @[AxiLoadQueue.scala 151:68:@13332.4]
  wire  _T_15386; // @[AxiLoadQueue.scala 150:92:@13334.4]
  wire  _T_15387; // @[AxiLoadQueue.scala 151:41:@13335.4]
  wire  _T_15388; // @[AxiLoadQueue.scala 152:30:@13336.4]
  wire  conflict_13_1; // @[AxiLoadQueue.scala 151:68:@13337.4]
  wire  _T_15390; // @[AxiLoadQueue.scala 150:92:@13339.4]
  wire  _T_15391; // @[AxiLoadQueue.scala 151:41:@13340.4]
  wire  _T_15392; // @[AxiLoadQueue.scala 152:30:@13341.4]
  wire  conflict_13_2; // @[AxiLoadQueue.scala 151:68:@13342.4]
  wire  _T_15394; // @[AxiLoadQueue.scala 150:92:@13344.4]
  wire  _T_15395; // @[AxiLoadQueue.scala 151:41:@13345.4]
  wire  _T_15396; // @[AxiLoadQueue.scala 152:30:@13346.4]
  wire  conflict_13_3; // @[AxiLoadQueue.scala 151:68:@13347.4]
  wire  _T_15398; // @[AxiLoadQueue.scala 150:92:@13349.4]
  wire  _T_15399; // @[AxiLoadQueue.scala 151:41:@13350.4]
  wire  _T_15400; // @[AxiLoadQueue.scala 152:30:@13351.4]
  wire  conflict_13_4; // @[AxiLoadQueue.scala 151:68:@13352.4]
  wire  _T_15402; // @[AxiLoadQueue.scala 150:92:@13354.4]
  wire  _T_15403; // @[AxiLoadQueue.scala 151:41:@13355.4]
  wire  _T_15404; // @[AxiLoadQueue.scala 152:30:@13356.4]
  wire  conflict_13_5; // @[AxiLoadQueue.scala 151:68:@13357.4]
  wire  _T_15406; // @[AxiLoadQueue.scala 150:92:@13359.4]
  wire  _T_15407; // @[AxiLoadQueue.scala 151:41:@13360.4]
  wire  _T_15408; // @[AxiLoadQueue.scala 152:30:@13361.4]
  wire  conflict_13_6; // @[AxiLoadQueue.scala 151:68:@13362.4]
  wire  _T_15410; // @[AxiLoadQueue.scala 150:92:@13364.4]
  wire  _T_15411; // @[AxiLoadQueue.scala 151:41:@13365.4]
  wire  _T_15412; // @[AxiLoadQueue.scala 152:30:@13366.4]
  wire  conflict_13_7; // @[AxiLoadQueue.scala 151:68:@13367.4]
  wire  _T_15414; // @[AxiLoadQueue.scala 150:92:@13369.4]
  wire  _T_15415; // @[AxiLoadQueue.scala 151:41:@13370.4]
  wire  _T_15416; // @[AxiLoadQueue.scala 152:30:@13371.4]
  wire  conflict_13_8; // @[AxiLoadQueue.scala 151:68:@13372.4]
  wire  _T_15418; // @[AxiLoadQueue.scala 150:92:@13374.4]
  wire  _T_15419; // @[AxiLoadQueue.scala 151:41:@13375.4]
  wire  _T_15420; // @[AxiLoadQueue.scala 152:30:@13376.4]
  wire  conflict_13_9; // @[AxiLoadQueue.scala 151:68:@13377.4]
  wire  _T_15422; // @[AxiLoadQueue.scala 150:92:@13379.4]
  wire  _T_15423; // @[AxiLoadQueue.scala 151:41:@13380.4]
  wire  _T_15424; // @[AxiLoadQueue.scala 152:30:@13381.4]
  wire  conflict_13_10; // @[AxiLoadQueue.scala 151:68:@13382.4]
  wire  _T_15426; // @[AxiLoadQueue.scala 150:92:@13384.4]
  wire  _T_15427; // @[AxiLoadQueue.scala 151:41:@13385.4]
  wire  _T_15428; // @[AxiLoadQueue.scala 152:30:@13386.4]
  wire  conflict_13_11; // @[AxiLoadQueue.scala 151:68:@13387.4]
  wire  _T_15430; // @[AxiLoadQueue.scala 150:92:@13389.4]
  wire  _T_15431; // @[AxiLoadQueue.scala 151:41:@13390.4]
  wire  _T_15432; // @[AxiLoadQueue.scala 152:30:@13391.4]
  wire  conflict_13_12; // @[AxiLoadQueue.scala 151:68:@13392.4]
  wire  _T_15434; // @[AxiLoadQueue.scala 150:92:@13394.4]
  wire  _T_15435; // @[AxiLoadQueue.scala 151:41:@13395.4]
  wire  _T_15436; // @[AxiLoadQueue.scala 152:30:@13396.4]
  wire  conflict_13_13; // @[AxiLoadQueue.scala 151:68:@13397.4]
  wire  _T_15438; // @[AxiLoadQueue.scala 150:92:@13399.4]
  wire  _T_15439; // @[AxiLoadQueue.scala 151:41:@13400.4]
  wire  _T_15440; // @[AxiLoadQueue.scala 152:30:@13401.4]
  wire  conflict_13_14; // @[AxiLoadQueue.scala 151:68:@13402.4]
  wire  _T_15442; // @[AxiLoadQueue.scala 150:92:@13404.4]
  wire  _T_15443; // @[AxiLoadQueue.scala 151:41:@13405.4]
  wire  _T_15444; // @[AxiLoadQueue.scala 152:30:@13406.4]
  wire  conflict_13_15; // @[AxiLoadQueue.scala 151:68:@13407.4]
  wire  _T_15446; // @[AxiLoadQueue.scala 150:92:@13409.4]
  wire  _T_15447; // @[AxiLoadQueue.scala 151:41:@13410.4]
  wire  _T_15448; // @[AxiLoadQueue.scala 152:30:@13411.4]
  wire  conflict_14_0; // @[AxiLoadQueue.scala 151:68:@13412.4]
  wire  _T_15450; // @[AxiLoadQueue.scala 150:92:@13414.4]
  wire  _T_15451; // @[AxiLoadQueue.scala 151:41:@13415.4]
  wire  _T_15452; // @[AxiLoadQueue.scala 152:30:@13416.4]
  wire  conflict_14_1; // @[AxiLoadQueue.scala 151:68:@13417.4]
  wire  _T_15454; // @[AxiLoadQueue.scala 150:92:@13419.4]
  wire  _T_15455; // @[AxiLoadQueue.scala 151:41:@13420.4]
  wire  _T_15456; // @[AxiLoadQueue.scala 152:30:@13421.4]
  wire  conflict_14_2; // @[AxiLoadQueue.scala 151:68:@13422.4]
  wire  _T_15458; // @[AxiLoadQueue.scala 150:92:@13424.4]
  wire  _T_15459; // @[AxiLoadQueue.scala 151:41:@13425.4]
  wire  _T_15460; // @[AxiLoadQueue.scala 152:30:@13426.4]
  wire  conflict_14_3; // @[AxiLoadQueue.scala 151:68:@13427.4]
  wire  _T_15462; // @[AxiLoadQueue.scala 150:92:@13429.4]
  wire  _T_15463; // @[AxiLoadQueue.scala 151:41:@13430.4]
  wire  _T_15464; // @[AxiLoadQueue.scala 152:30:@13431.4]
  wire  conflict_14_4; // @[AxiLoadQueue.scala 151:68:@13432.4]
  wire  _T_15466; // @[AxiLoadQueue.scala 150:92:@13434.4]
  wire  _T_15467; // @[AxiLoadQueue.scala 151:41:@13435.4]
  wire  _T_15468; // @[AxiLoadQueue.scala 152:30:@13436.4]
  wire  conflict_14_5; // @[AxiLoadQueue.scala 151:68:@13437.4]
  wire  _T_15470; // @[AxiLoadQueue.scala 150:92:@13439.4]
  wire  _T_15471; // @[AxiLoadQueue.scala 151:41:@13440.4]
  wire  _T_15472; // @[AxiLoadQueue.scala 152:30:@13441.4]
  wire  conflict_14_6; // @[AxiLoadQueue.scala 151:68:@13442.4]
  wire  _T_15474; // @[AxiLoadQueue.scala 150:92:@13444.4]
  wire  _T_15475; // @[AxiLoadQueue.scala 151:41:@13445.4]
  wire  _T_15476; // @[AxiLoadQueue.scala 152:30:@13446.4]
  wire  conflict_14_7; // @[AxiLoadQueue.scala 151:68:@13447.4]
  wire  _T_15478; // @[AxiLoadQueue.scala 150:92:@13449.4]
  wire  _T_15479; // @[AxiLoadQueue.scala 151:41:@13450.4]
  wire  _T_15480; // @[AxiLoadQueue.scala 152:30:@13451.4]
  wire  conflict_14_8; // @[AxiLoadQueue.scala 151:68:@13452.4]
  wire  _T_15482; // @[AxiLoadQueue.scala 150:92:@13454.4]
  wire  _T_15483; // @[AxiLoadQueue.scala 151:41:@13455.4]
  wire  _T_15484; // @[AxiLoadQueue.scala 152:30:@13456.4]
  wire  conflict_14_9; // @[AxiLoadQueue.scala 151:68:@13457.4]
  wire  _T_15486; // @[AxiLoadQueue.scala 150:92:@13459.4]
  wire  _T_15487; // @[AxiLoadQueue.scala 151:41:@13460.4]
  wire  _T_15488; // @[AxiLoadQueue.scala 152:30:@13461.4]
  wire  conflict_14_10; // @[AxiLoadQueue.scala 151:68:@13462.4]
  wire  _T_15490; // @[AxiLoadQueue.scala 150:92:@13464.4]
  wire  _T_15491; // @[AxiLoadQueue.scala 151:41:@13465.4]
  wire  _T_15492; // @[AxiLoadQueue.scala 152:30:@13466.4]
  wire  conflict_14_11; // @[AxiLoadQueue.scala 151:68:@13467.4]
  wire  _T_15494; // @[AxiLoadQueue.scala 150:92:@13469.4]
  wire  _T_15495; // @[AxiLoadQueue.scala 151:41:@13470.4]
  wire  _T_15496; // @[AxiLoadQueue.scala 152:30:@13471.4]
  wire  conflict_14_12; // @[AxiLoadQueue.scala 151:68:@13472.4]
  wire  _T_15498; // @[AxiLoadQueue.scala 150:92:@13474.4]
  wire  _T_15499; // @[AxiLoadQueue.scala 151:41:@13475.4]
  wire  _T_15500; // @[AxiLoadQueue.scala 152:30:@13476.4]
  wire  conflict_14_13; // @[AxiLoadQueue.scala 151:68:@13477.4]
  wire  _T_15502; // @[AxiLoadQueue.scala 150:92:@13479.4]
  wire  _T_15503; // @[AxiLoadQueue.scala 151:41:@13480.4]
  wire  _T_15504; // @[AxiLoadQueue.scala 152:30:@13481.4]
  wire  conflict_14_14; // @[AxiLoadQueue.scala 151:68:@13482.4]
  wire  _T_15506; // @[AxiLoadQueue.scala 150:92:@13484.4]
  wire  _T_15507; // @[AxiLoadQueue.scala 151:41:@13485.4]
  wire  _T_15508; // @[AxiLoadQueue.scala 152:30:@13486.4]
  wire  conflict_14_15; // @[AxiLoadQueue.scala 151:68:@13487.4]
  wire  _T_15510; // @[AxiLoadQueue.scala 150:92:@13489.4]
  wire  _T_15511; // @[AxiLoadQueue.scala 151:41:@13490.4]
  wire  _T_15512; // @[AxiLoadQueue.scala 152:30:@13491.4]
  wire  conflict_15_0; // @[AxiLoadQueue.scala 151:68:@13492.4]
  wire  _T_15514; // @[AxiLoadQueue.scala 150:92:@13494.4]
  wire  _T_15515; // @[AxiLoadQueue.scala 151:41:@13495.4]
  wire  _T_15516; // @[AxiLoadQueue.scala 152:30:@13496.4]
  wire  conflict_15_1; // @[AxiLoadQueue.scala 151:68:@13497.4]
  wire  _T_15518; // @[AxiLoadQueue.scala 150:92:@13499.4]
  wire  _T_15519; // @[AxiLoadQueue.scala 151:41:@13500.4]
  wire  _T_15520; // @[AxiLoadQueue.scala 152:30:@13501.4]
  wire  conflict_15_2; // @[AxiLoadQueue.scala 151:68:@13502.4]
  wire  _T_15522; // @[AxiLoadQueue.scala 150:92:@13504.4]
  wire  _T_15523; // @[AxiLoadQueue.scala 151:41:@13505.4]
  wire  _T_15524; // @[AxiLoadQueue.scala 152:30:@13506.4]
  wire  conflict_15_3; // @[AxiLoadQueue.scala 151:68:@13507.4]
  wire  _T_15526; // @[AxiLoadQueue.scala 150:92:@13509.4]
  wire  _T_15527; // @[AxiLoadQueue.scala 151:41:@13510.4]
  wire  _T_15528; // @[AxiLoadQueue.scala 152:30:@13511.4]
  wire  conflict_15_4; // @[AxiLoadQueue.scala 151:68:@13512.4]
  wire  _T_15530; // @[AxiLoadQueue.scala 150:92:@13514.4]
  wire  _T_15531; // @[AxiLoadQueue.scala 151:41:@13515.4]
  wire  _T_15532; // @[AxiLoadQueue.scala 152:30:@13516.4]
  wire  conflict_15_5; // @[AxiLoadQueue.scala 151:68:@13517.4]
  wire  _T_15534; // @[AxiLoadQueue.scala 150:92:@13519.4]
  wire  _T_15535; // @[AxiLoadQueue.scala 151:41:@13520.4]
  wire  _T_15536; // @[AxiLoadQueue.scala 152:30:@13521.4]
  wire  conflict_15_6; // @[AxiLoadQueue.scala 151:68:@13522.4]
  wire  _T_15538; // @[AxiLoadQueue.scala 150:92:@13524.4]
  wire  _T_15539; // @[AxiLoadQueue.scala 151:41:@13525.4]
  wire  _T_15540; // @[AxiLoadQueue.scala 152:30:@13526.4]
  wire  conflict_15_7; // @[AxiLoadQueue.scala 151:68:@13527.4]
  wire  _T_15542; // @[AxiLoadQueue.scala 150:92:@13529.4]
  wire  _T_15543; // @[AxiLoadQueue.scala 151:41:@13530.4]
  wire  _T_15544; // @[AxiLoadQueue.scala 152:30:@13531.4]
  wire  conflict_15_8; // @[AxiLoadQueue.scala 151:68:@13532.4]
  wire  _T_15546; // @[AxiLoadQueue.scala 150:92:@13534.4]
  wire  _T_15547; // @[AxiLoadQueue.scala 151:41:@13535.4]
  wire  _T_15548; // @[AxiLoadQueue.scala 152:30:@13536.4]
  wire  conflict_15_9; // @[AxiLoadQueue.scala 151:68:@13537.4]
  wire  _T_15550; // @[AxiLoadQueue.scala 150:92:@13539.4]
  wire  _T_15551; // @[AxiLoadQueue.scala 151:41:@13540.4]
  wire  _T_15552; // @[AxiLoadQueue.scala 152:30:@13541.4]
  wire  conflict_15_10; // @[AxiLoadQueue.scala 151:68:@13542.4]
  wire  _T_15554; // @[AxiLoadQueue.scala 150:92:@13544.4]
  wire  _T_15555; // @[AxiLoadQueue.scala 151:41:@13545.4]
  wire  _T_15556; // @[AxiLoadQueue.scala 152:30:@13546.4]
  wire  conflict_15_11; // @[AxiLoadQueue.scala 151:68:@13547.4]
  wire  _T_15558; // @[AxiLoadQueue.scala 150:92:@13549.4]
  wire  _T_15559; // @[AxiLoadQueue.scala 151:41:@13550.4]
  wire  _T_15560; // @[AxiLoadQueue.scala 152:30:@13551.4]
  wire  conflict_15_12; // @[AxiLoadQueue.scala 151:68:@13552.4]
  wire  _T_15562; // @[AxiLoadQueue.scala 150:92:@13554.4]
  wire  _T_15563; // @[AxiLoadQueue.scala 151:41:@13555.4]
  wire  _T_15564; // @[AxiLoadQueue.scala 152:30:@13556.4]
  wire  conflict_15_13; // @[AxiLoadQueue.scala 151:68:@13557.4]
  wire  _T_15566; // @[AxiLoadQueue.scala 150:92:@13559.4]
  wire  _T_15567; // @[AxiLoadQueue.scala 151:41:@13560.4]
  wire  _T_15568; // @[AxiLoadQueue.scala 152:30:@13561.4]
  wire  conflict_15_14; // @[AxiLoadQueue.scala 151:68:@13562.4]
  wire  _T_15570; // @[AxiLoadQueue.scala 150:92:@13564.4]
  wire  _T_15571; // @[AxiLoadQueue.scala 151:41:@13565.4]
  wire  _T_15572; // @[AxiLoadQueue.scala 152:30:@13566.4]
  wire  conflict_15_15; // @[AxiLoadQueue.scala 151:68:@13567.4]
  wire  _T_16805; // @[AxiLoadQueue.scala 163:13:@13570.4]
  wire  storeAddrNotKnownFlags_0_0; // @[AxiLoadQueue.scala 163:19:@13571.4]
  wire  _T_16808; // @[AxiLoadQueue.scala 163:13:@13572.4]
  wire  storeAddrNotKnownFlags_0_1; // @[AxiLoadQueue.scala 163:19:@13573.4]
  wire  _T_16811; // @[AxiLoadQueue.scala 163:13:@13574.4]
  wire  storeAddrNotKnownFlags_0_2; // @[AxiLoadQueue.scala 163:19:@13575.4]
  wire  _T_16814; // @[AxiLoadQueue.scala 163:13:@13576.4]
  wire  storeAddrNotKnownFlags_0_3; // @[AxiLoadQueue.scala 163:19:@13577.4]
  wire  _T_16817; // @[AxiLoadQueue.scala 163:13:@13578.4]
  wire  storeAddrNotKnownFlags_0_4; // @[AxiLoadQueue.scala 163:19:@13579.4]
  wire  _T_16820; // @[AxiLoadQueue.scala 163:13:@13580.4]
  wire  storeAddrNotKnownFlags_0_5; // @[AxiLoadQueue.scala 163:19:@13581.4]
  wire  _T_16823; // @[AxiLoadQueue.scala 163:13:@13582.4]
  wire  storeAddrNotKnownFlags_0_6; // @[AxiLoadQueue.scala 163:19:@13583.4]
  wire  _T_16826; // @[AxiLoadQueue.scala 163:13:@13584.4]
  wire  storeAddrNotKnownFlags_0_7; // @[AxiLoadQueue.scala 163:19:@13585.4]
  wire  _T_16829; // @[AxiLoadQueue.scala 163:13:@13586.4]
  wire  storeAddrNotKnownFlags_0_8; // @[AxiLoadQueue.scala 163:19:@13587.4]
  wire  _T_16832; // @[AxiLoadQueue.scala 163:13:@13588.4]
  wire  storeAddrNotKnownFlags_0_9; // @[AxiLoadQueue.scala 163:19:@13589.4]
  wire  _T_16835; // @[AxiLoadQueue.scala 163:13:@13590.4]
  wire  storeAddrNotKnownFlags_0_10; // @[AxiLoadQueue.scala 163:19:@13591.4]
  wire  _T_16838; // @[AxiLoadQueue.scala 163:13:@13592.4]
  wire  storeAddrNotKnownFlags_0_11; // @[AxiLoadQueue.scala 163:19:@13593.4]
  wire  _T_16841; // @[AxiLoadQueue.scala 163:13:@13594.4]
  wire  storeAddrNotKnownFlags_0_12; // @[AxiLoadQueue.scala 163:19:@13595.4]
  wire  _T_16844; // @[AxiLoadQueue.scala 163:13:@13596.4]
  wire  storeAddrNotKnownFlags_0_13; // @[AxiLoadQueue.scala 163:19:@13597.4]
  wire  _T_16847; // @[AxiLoadQueue.scala 163:13:@13598.4]
  wire  storeAddrNotKnownFlags_0_14; // @[AxiLoadQueue.scala 163:19:@13599.4]
  wire  _T_16850; // @[AxiLoadQueue.scala 163:13:@13600.4]
  wire  storeAddrNotKnownFlags_0_15; // @[AxiLoadQueue.scala 163:19:@13601.4]
  wire  storeAddrNotKnownFlags_1_0; // @[AxiLoadQueue.scala 163:19:@13619.4]
  wire  storeAddrNotKnownFlags_1_1; // @[AxiLoadQueue.scala 163:19:@13621.4]
  wire  storeAddrNotKnownFlags_1_2; // @[AxiLoadQueue.scala 163:19:@13623.4]
  wire  storeAddrNotKnownFlags_1_3; // @[AxiLoadQueue.scala 163:19:@13625.4]
  wire  storeAddrNotKnownFlags_1_4; // @[AxiLoadQueue.scala 163:19:@13627.4]
  wire  storeAddrNotKnownFlags_1_5; // @[AxiLoadQueue.scala 163:19:@13629.4]
  wire  storeAddrNotKnownFlags_1_6; // @[AxiLoadQueue.scala 163:19:@13631.4]
  wire  storeAddrNotKnownFlags_1_7; // @[AxiLoadQueue.scala 163:19:@13633.4]
  wire  storeAddrNotKnownFlags_1_8; // @[AxiLoadQueue.scala 163:19:@13635.4]
  wire  storeAddrNotKnownFlags_1_9; // @[AxiLoadQueue.scala 163:19:@13637.4]
  wire  storeAddrNotKnownFlags_1_10; // @[AxiLoadQueue.scala 163:19:@13639.4]
  wire  storeAddrNotKnownFlags_1_11; // @[AxiLoadQueue.scala 163:19:@13641.4]
  wire  storeAddrNotKnownFlags_1_12; // @[AxiLoadQueue.scala 163:19:@13643.4]
  wire  storeAddrNotKnownFlags_1_13; // @[AxiLoadQueue.scala 163:19:@13645.4]
  wire  storeAddrNotKnownFlags_1_14; // @[AxiLoadQueue.scala 163:19:@13647.4]
  wire  storeAddrNotKnownFlags_1_15; // @[AxiLoadQueue.scala 163:19:@13649.4]
  wire  storeAddrNotKnownFlags_2_0; // @[AxiLoadQueue.scala 163:19:@13667.4]
  wire  storeAddrNotKnownFlags_2_1; // @[AxiLoadQueue.scala 163:19:@13669.4]
  wire  storeAddrNotKnownFlags_2_2; // @[AxiLoadQueue.scala 163:19:@13671.4]
  wire  storeAddrNotKnownFlags_2_3; // @[AxiLoadQueue.scala 163:19:@13673.4]
  wire  storeAddrNotKnownFlags_2_4; // @[AxiLoadQueue.scala 163:19:@13675.4]
  wire  storeAddrNotKnownFlags_2_5; // @[AxiLoadQueue.scala 163:19:@13677.4]
  wire  storeAddrNotKnownFlags_2_6; // @[AxiLoadQueue.scala 163:19:@13679.4]
  wire  storeAddrNotKnownFlags_2_7; // @[AxiLoadQueue.scala 163:19:@13681.4]
  wire  storeAddrNotKnownFlags_2_8; // @[AxiLoadQueue.scala 163:19:@13683.4]
  wire  storeAddrNotKnownFlags_2_9; // @[AxiLoadQueue.scala 163:19:@13685.4]
  wire  storeAddrNotKnownFlags_2_10; // @[AxiLoadQueue.scala 163:19:@13687.4]
  wire  storeAddrNotKnownFlags_2_11; // @[AxiLoadQueue.scala 163:19:@13689.4]
  wire  storeAddrNotKnownFlags_2_12; // @[AxiLoadQueue.scala 163:19:@13691.4]
  wire  storeAddrNotKnownFlags_2_13; // @[AxiLoadQueue.scala 163:19:@13693.4]
  wire  storeAddrNotKnownFlags_2_14; // @[AxiLoadQueue.scala 163:19:@13695.4]
  wire  storeAddrNotKnownFlags_2_15; // @[AxiLoadQueue.scala 163:19:@13697.4]
  wire  storeAddrNotKnownFlags_3_0; // @[AxiLoadQueue.scala 163:19:@13715.4]
  wire  storeAddrNotKnownFlags_3_1; // @[AxiLoadQueue.scala 163:19:@13717.4]
  wire  storeAddrNotKnownFlags_3_2; // @[AxiLoadQueue.scala 163:19:@13719.4]
  wire  storeAddrNotKnownFlags_3_3; // @[AxiLoadQueue.scala 163:19:@13721.4]
  wire  storeAddrNotKnownFlags_3_4; // @[AxiLoadQueue.scala 163:19:@13723.4]
  wire  storeAddrNotKnownFlags_3_5; // @[AxiLoadQueue.scala 163:19:@13725.4]
  wire  storeAddrNotKnownFlags_3_6; // @[AxiLoadQueue.scala 163:19:@13727.4]
  wire  storeAddrNotKnownFlags_3_7; // @[AxiLoadQueue.scala 163:19:@13729.4]
  wire  storeAddrNotKnownFlags_3_8; // @[AxiLoadQueue.scala 163:19:@13731.4]
  wire  storeAddrNotKnownFlags_3_9; // @[AxiLoadQueue.scala 163:19:@13733.4]
  wire  storeAddrNotKnownFlags_3_10; // @[AxiLoadQueue.scala 163:19:@13735.4]
  wire  storeAddrNotKnownFlags_3_11; // @[AxiLoadQueue.scala 163:19:@13737.4]
  wire  storeAddrNotKnownFlags_3_12; // @[AxiLoadQueue.scala 163:19:@13739.4]
  wire  storeAddrNotKnownFlags_3_13; // @[AxiLoadQueue.scala 163:19:@13741.4]
  wire  storeAddrNotKnownFlags_3_14; // @[AxiLoadQueue.scala 163:19:@13743.4]
  wire  storeAddrNotKnownFlags_3_15; // @[AxiLoadQueue.scala 163:19:@13745.4]
  wire  storeAddrNotKnownFlags_4_0; // @[AxiLoadQueue.scala 163:19:@13763.4]
  wire  storeAddrNotKnownFlags_4_1; // @[AxiLoadQueue.scala 163:19:@13765.4]
  wire  storeAddrNotKnownFlags_4_2; // @[AxiLoadQueue.scala 163:19:@13767.4]
  wire  storeAddrNotKnownFlags_4_3; // @[AxiLoadQueue.scala 163:19:@13769.4]
  wire  storeAddrNotKnownFlags_4_4; // @[AxiLoadQueue.scala 163:19:@13771.4]
  wire  storeAddrNotKnownFlags_4_5; // @[AxiLoadQueue.scala 163:19:@13773.4]
  wire  storeAddrNotKnownFlags_4_6; // @[AxiLoadQueue.scala 163:19:@13775.4]
  wire  storeAddrNotKnownFlags_4_7; // @[AxiLoadQueue.scala 163:19:@13777.4]
  wire  storeAddrNotKnownFlags_4_8; // @[AxiLoadQueue.scala 163:19:@13779.4]
  wire  storeAddrNotKnownFlags_4_9; // @[AxiLoadQueue.scala 163:19:@13781.4]
  wire  storeAddrNotKnownFlags_4_10; // @[AxiLoadQueue.scala 163:19:@13783.4]
  wire  storeAddrNotKnownFlags_4_11; // @[AxiLoadQueue.scala 163:19:@13785.4]
  wire  storeAddrNotKnownFlags_4_12; // @[AxiLoadQueue.scala 163:19:@13787.4]
  wire  storeAddrNotKnownFlags_4_13; // @[AxiLoadQueue.scala 163:19:@13789.4]
  wire  storeAddrNotKnownFlags_4_14; // @[AxiLoadQueue.scala 163:19:@13791.4]
  wire  storeAddrNotKnownFlags_4_15; // @[AxiLoadQueue.scala 163:19:@13793.4]
  wire  storeAddrNotKnownFlags_5_0; // @[AxiLoadQueue.scala 163:19:@13811.4]
  wire  storeAddrNotKnownFlags_5_1; // @[AxiLoadQueue.scala 163:19:@13813.4]
  wire  storeAddrNotKnownFlags_5_2; // @[AxiLoadQueue.scala 163:19:@13815.4]
  wire  storeAddrNotKnownFlags_5_3; // @[AxiLoadQueue.scala 163:19:@13817.4]
  wire  storeAddrNotKnownFlags_5_4; // @[AxiLoadQueue.scala 163:19:@13819.4]
  wire  storeAddrNotKnownFlags_5_5; // @[AxiLoadQueue.scala 163:19:@13821.4]
  wire  storeAddrNotKnownFlags_5_6; // @[AxiLoadQueue.scala 163:19:@13823.4]
  wire  storeAddrNotKnownFlags_5_7; // @[AxiLoadQueue.scala 163:19:@13825.4]
  wire  storeAddrNotKnownFlags_5_8; // @[AxiLoadQueue.scala 163:19:@13827.4]
  wire  storeAddrNotKnownFlags_5_9; // @[AxiLoadQueue.scala 163:19:@13829.4]
  wire  storeAddrNotKnownFlags_5_10; // @[AxiLoadQueue.scala 163:19:@13831.4]
  wire  storeAddrNotKnownFlags_5_11; // @[AxiLoadQueue.scala 163:19:@13833.4]
  wire  storeAddrNotKnownFlags_5_12; // @[AxiLoadQueue.scala 163:19:@13835.4]
  wire  storeAddrNotKnownFlags_5_13; // @[AxiLoadQueue.scala 163:19:@13837.4]
  wire  storeAddrNotKnownFlags_5_14; // @[AxiLoadQueue.scala 163:19:@13839.4]
  wire  storeAddrNotKnownFlags_5_15; // @[AxiLoadQueue.scala 163:19:@13841.4]
  wire  storeAddrNotKnownFlags_6_0; // @[AxiLoadQueue.scala 163:19:@13859.4]
  wire  storeAddrNotKnownFlags_6_1; // @[AxiLoadQueue.scala 163:19:@13861.4]
  wire  storeAddrNotKnownFlags_6_2; // @[AxiLoadQueue.scala 163:19:@13863.4]
  wire  storeAddrNotKnownFlags_6_3; // @[AxiLoadQueue.scala 163:19:@13865.4]
  wire  storeAddrNotKnownFlags_6_4; // @[AxiLoadQueue.scala 163:19:@13867.4]
  wire  storeAddrNotKnownFlags_6_5; // @[AxiLoadQueue.scala 163:19:@13869.4]
  wire  storeAddrNotKnownFlags_6_6; // @[AxiLoadQueue.scala 163:19:@13871.4]
  wire  storeAddrNotKnownFlags_6_7; // @[AxiLoadQueue.scala 163:19:@13873.4]
  wire  storeAddrNotKnownFlags_6_8; // @[AxiLoadQueue.scala 163:19:@13875.4]
  wire  storeAddrNotKnownFlags_6_9; // @[AxiLoadQueue.scala 163:19:@13877.4]
  wire  storeAddrNotKnownFlags_6_10; // @[AxiLoadQueue.scala 163:19:@13879.4]
  wire  storeAddrNotKnownFlags_6_11; // @[AxiLoadQueue.scala 163:19:@13881.4]
  wire  storeAddrNotKnownFlags_6_12; // @[AxiLoadQueue.scala 163:19:@13883.4]
  wire  storeAddrNotKnownFlags_6_13; // @[AxiLoadQueue.scala 163:19:@13885.4]
  wire  storeAddrNotKnownFlags_6_14; // @[AxiLoadQueue.scala 163:19:@13887.4]
  wire  storeAddrNotKnownFlags_6_15; // @[AxiLoadQueue.scala 163:19:@13889.4]
  wire  storeAddrNotKnownFlags_7_0; // @[AxiLoadQueue.scala 163:19:@13907.4]
  wire  storeAddrNotKnownFlags_7_1; // @[AxiLoadQueue.scala 163:19:@13909.4]
  wire  storeAddrNotKnownFlags_7_2; // @[AxiLoadQueue.scala 163:19:@13911.4]
  wire  storeAddrNotKnownFlags_7_3; // @[AxiLoadQueue.scala 163:19:@13913.4]
  wire  storeAddrNotKnownFlags_7_4; // @[AxiLoadQueue.scala 163:19:@13915.4]
  wire  storeAddrNotKnownFlags_7_5; // @[AxiLoadQueue.scala 163:19:@13917.4]
  wire  storeAddrNotKnownFlags_7_6; // @[AxiLoadQueue.scala 163:19:@13919.4]
  wire  storeAddrNotKnownFlags_7_7; // @[AxiLoadQueue.scala 163:19:@13921.4]
  wire  storeAddrNotKnownFlags_7_8; // @[AxiLoadQueue.scala 163:19:@13923.4]
  wire  storeAddrNotKnownFlags_7_9; // @[AxiLoadQueue.scala 163:19:@13925.4]
  wire  storeAddrNotKnownFlags_7_10; // @[AxiLoadQueue.scala 163:19:@13927.4]
  wire  storeAddrNotKnownFlags_7_11; // @[AxiLoadQueue.scala 163:19:@13929.4]
  wire  storeAddrNotKnownFlags_7_12; // @[AxiLoadQueue.scala 163:19:@13931.4]
  wire  storeAddrNotKnownFlags_7_13; // @[AxiLoadQueue.scala 163:19:@13933.4]
  wire  storeAddrNotKnownFlags_7_14; // @[AxiLoadQueue.scala 163:19:@13935.4]
  wire  storeAddrNotKnownFlags_7_15; // @[AxiLoadQueue.scala 163:19:@13937.4]
  wire  storeAddrNotKnownFlags_8_0; // @[AxiLoadQueue.scala 163:19:@13955.4]
  wire  storeAddrNotKnownFlags_8_1; // @[AxiLoadQueue.scala 163:19:@13957.4]
  wire  storeAddrNotKnownFlags_8_2; // @[AxiLoadQueue.scala 163:19:@13959.4]
  wire  storeAddrNotKnownFlags_8_3; // @[AxiLoadQueue.scala 163:19:@13961.4]
  wire  storeAddrNotKnownFlags_8_4; // @[AxiLoadQueue.scala 163:19:@13963.4]
  wire  storeAddrNotKnownFlags_8_5; // @[AxiLoadQueue.scala 163:19:@13965.4]
  wire  storeAddrNotKnownFlags_8_6; // @[AxiLoadQueue.scala 163:19:@13967.4]
  wire  storeAddrNotKnownFlags_8_7; // @[AxiLoadQueue.scala 163:19:@13969.4]
  wire  storeAddrNotKnownFlags_8_8; // @[AxiLoadQueue.scala 163:19:@13971.4]
  wire  storeAddrNotKnownFlags_8_9; // @[AxiLoadQueue.scala 163:19:@13973.4]
  wire  storeAddrNotKnownFlags_8_10; // @[AxiLoadQueue.scala 163:19:@13975.4]
  wire  storeAddrNotKnownFlags_8_11; // @[AxiLoadQueue.scala 163:19:@13977.4]
  wire  storeAddrNotKnownFlags_8_12; // @[AxiLoadQueue.scala 163:19:@13979.4]
  wire  storeAddrNotKnownFlags_8_13; // @[AxiLoadQueue.scala 163:19:@13981.4]
  wire  storeAddrNotKnownFlags_8_14; // @[AxiLoadQueue.scala 163:19:@13983.4]
  wire  storeAddrNotKnownFlags_8_15; // @[AxiLoadQueue.scala 163:19:@13985.4]
  wire  storeAddrNotKnownFlags_9_0; // @[AxiLoadQueue.scala 163:19:@14003.4]
  wire  storeAddrNotKnownFlags_9_1; // @[AxiLoadQueue.scala 163:19:@14005.4]
  wire  storeAddrNotKnownFlags_9_2; // @[AxiLoadQueue.scala 163:19:@14007.4]
  wire  storeAddrNotKnownFlags_9_3; // @[AxiLoadQueue.scala 163:19:@14009.4]
  wire  storeAddrNotKnownFlags_9_4; // @[AxiLoadQueue.scala 163:19:@14011.4]
  wire  storeAddrNotKnownFlags_9_5; // @[AxiLoadQueue.scala 163:19:@14013.4]
  wire  storeAddrNotKnownFlags_9_6; // @[AxiLoadQueue.scala 163:19:@14015.4]
  wire  storeAddrNotKnownFlags_9_7; // @[AxiLoadQueue.scala 163:19:@14017.4]
  wire  storeAddrNotKnownFlags_9_8; // @[AxiLoadQueue.scala 163:19:@14019.4]
  wire  storeAddrNotKnownFlags_9_9; // @[AxiLoadQueue.scala 163:19:@14021.4]
  wire  storeAddrNotKnownFlags_9_10; // @[AxiLoadQueue.scala 163:19:@14023.4]
  wire  storeAddrNotKnownFlags_9_11; // @[AxiLoadQueue.scala 163:19:@14025.4]
  wire  storeAddrNotKnownFlags_9_12; // @[AxiLoadQueue.scala 163:19:@14027.4]
  wire  storeAddrNotKnownFlags_9_13; // @[AxiLoadQueue.scala 163:19:@14029.4]
  wire  storeAddrNotKnownFlags_9_14; // @[AxiLoadQueue.scala 163:19:@14031.4]
  wire  storeAddrNotKnownFlags_9_15; // @[AxiLoadQueue.scala 163:19:@14033.4]
  wire  storeAddrNotKnownFlags_10_0; // @[AxiLoadQueue.scala 163:19:@14051.4]
  wire  storeAddrNotKnownFlags_10_1; // @[AxiLoadQueue.scala 163:19:@14053.4]
  wire  storeAddrNotKnownFlags_10_2; // @[AxiLoadQueue.scala 163:19:@14055.4]
  wire  storeAddrNotKnownFlags_10_3; // @[AxiLoadQueue.scala 163:19:@14057.4]
  wire  storeAddrNotKnownFlags_10_4; // @[AxiLoadQueue.scala 163:19:@14059.4]
  wire  storeAddrNotKnownFlags_10_5; // @[AxiLoadQueue.scala 163:19:@14061.4]
  wire  storeAddrNotKnownFlags_10_6; // @[AxiLoadQueue.scala 163:19:@14063.4]
  wire  storeAddrNotKnownFlags_10_7; // @[AxiLoadQueue.scala 163:19:@14065.4]
  wire  storeAddrNotKnownFlags_10_8; // @[AxiLoadQueue.scala 163:19:@14067.4]
  wire  storeAddrNotKnownFlags_10_9; // @[AxiLoadQueue.scala 163:19:@14069.4]
  wire  storeAddrNotKnownFlags_10_10; // @[AxiLoadQueue.scala 163:19:@14071.4]
  wire  storeAddrNotKnownFlags_10_11; // @[AxiLoadQueue.scala 163:19:@14073.4]
  wire  storeAddrNotKnownFlags_10_12; // @[AxiLoadQueue.scala 163:19:@14075.4]
  wire  storeAddrNotKnownFlags_10_13; // @[AxiLoadQueue.scala 163:19:@14077.4]
  wire  storeAddrNotKnownFlags_10_14; // @[AxiLoadQueue.scala 163:19:@14079.4]
  wire  storeAddrNotKnownFlags_10_15; // @[AxiLoadQueue.scala 163:19:@14081.4]
  wire  storeAddrNotKnownFlags_11_0; // @[AxiLoadQueue.scala 163:19:@14099.4]
  wire  storeAddrNotKnownFlags_11_1; // @[AxiLoadQueue.scala 163:19:@14101.4]
  wire  storeAddrNotKnownFlags_11_2; // @[AxiLoadQueue.scala 163:19:@14103.4]
  wire  storeAddrNotKnownFlags_11_3; // @[AxiLoadQueue.scala 163:19:@14105.4]
  wire  storeAddrNotKnownFlags_11_4; // @[AxiLoadQueue.scala 163:19:@14107.4]
  wire  storeAddrNotKnownFlags_11_5; // @[AxiLoadQueue.scala 163:19:@14109.4]
  wire  storeAddrNotKnownFlags_11_6; // @[AxiLoadQueue.scala 163:19:@14111.4]
  wire  storeAddrNotKnownFlags_11_7; // @[AxiLoadQueue.scala 163:19:@14113.4]
  wire  storeAddrNotKnownFlags_11_8; // @[AxiLoadQueue.scala 163:19:@14115.4]
  wire  storeAddrNotKnownFlags_11_9; // @[AxiLoadQueue.scala 163:19:@14117.4]
  wire  storeAddrNotKnownFlags_11_10; // @[AxiLoadQueue.scala 163:19:@14119.4]
  wire  storeAddrNotKnownFlags_11_11; // @[AxiLoadQueue.scala 163:19:@14121.4]
  wire  storeAddrNotKnownFlags_11_12; // @[AxiLoadQueue.scala 163:19:@14123.4]
  wire  storeAddrNotKnownFlags_11_13; // @[AxiLoadQueue.scala 163:19:@14125.4]
  wire  storeAddrNotKnownFlags_11_14; // @[AxiLoadQueue.scala 163:19:@14127.4]
  wire  storeAddrNotKnownFlags_11_15; // @[AxiLoadQueue.scala 163:19:@14129.4]
  wire  storeAddrNotKnownFlags_12_0; // @[AxiLoadQueue.scala 163:19:@14147.4]
  wire  storeAddrNotKnownFlags_12_1; // @[AxiLoadQueue.scala 163:19:@14149.4]
  wire  storeAddrNotKnownFlags_12_2; // @[AxiLoadQueue.scala 163:19:@14151.4]
  wire  storeAddrNotKnownFlags_12_3; // @[AxiLoadQueue.scala 163:19:@14153.4]
  wire  storeAddrNotKnownFlags_12_4; // @[AxiLoadQueue.scala 163:19:@14155.4]
  wire  storeAddrNotKnownFlags_12_5; // @[AxiLoadQueue.scala 163:19:@14157.4]
  wire  storeAddrNotKnownFlags_12_6; // @[AxiLoadQueue.scala 163:19:@14159.4]
  wire  storeAddrNotKnownFlags_12_7; // @[AxiLoadQueue.scala 163:19:@14161.4]
  wire  storeAddrNotKnownFlags_12_8; // @[AxiLoadQueue.scala 163:19:@14163.4]
  wire  storeAddrNotKnownFlags_12_9; // @[AxiLoadQueue.scala 163:19:@14165.4]
  wire  storeAddrNotKnownFlags_12_10; // @[AxiLoadQueue.scala 163:19:@14167.4]
  wire  storeAddrNotKnownFlags_12_11; // @[AxiLoadQueue.scala 163:19:@14169.4]
  wire  storeAddrNotKnownFlags_12_12; // @[AxiLoadQueue.scala 163:19:@14171.4]
  wire  storeAddrNotKnownFlags_12_13; // @[AxiLoadQueue.scala 163:19:@14173.4]
  wire  storeAddrNotKnownFlags_12_14; // @[AxiLoadQueue.scala 163:19:@14175.4]
  wire  storeAddrNotKnownFlags_12_15; // @[AxiLoadQueue.scala 163:19:@14177.4]
  wire  storeAddrNotKnownFlags_13_0; // @[AxiLoadQueue.scala 163:19:@14195.4]
  wire  storeAddrNotKnownFlags_13_1; // @[AxiLoadQueue.scala 163:19:@14197.4]
  wire  storeAddrNotKnownFlags_13_2; // @[AxiLoadQueue.scala 163:19:@14199.4]
  wire  storeAddrNotKnownFlags_13_3; // @[AxiLoadQueue.scala 163:19:@14201.4]
  wire  storeAddrNotKnownFlags_13_4; // @[AxiLoadQueue.scala 163:19:@14203.4]
  wire  storeAddrNotKnownFlags_13_5; // @[AxiLoadQueue.scala 163:19:@14205.4]
  wire  storeAddrNotKnownFlags_13_6; // @[AxiLoadQueue.scala 163:19:@14207.4]
  wire  storeAddrNotKnownFlags_13_7; // @[AxiLoadQueue.scala 163:19:@14209.4]
  wire  storeAddrNotKnownFlags_13_8; // @[AxiLoadQueue.scala 163:19:@14211.4]
  wire  storeAddrNotKnownFlags_13_9; // @[AxiLoadQueue.scala 163:19:@14213.4]
  wire  storeAddrNotKnownFlags_13_10; // @[AxiLoadQueue.scala 163:19:@14215.4]
  wire  storeAddrNotKnownFlags_13_11; // @[AxiLoadQueue.scala 163:19:@14217.4]
  wire  storeAddrNotKnownFlags_13_12; // @[AxiLoadQueue.scala 163:19:@14219.4]
  wire  storeAddrNotKnownFlags_13_13; // @[AxiLoadQueue.scala 163:19:@14221.4]
  wire  storeAddrNotKnownFlags_13_14; // @[AxiLoadQueue.scala 163:19:@14223.4]
  wire  storeAddrNotKnownFlags_13_15; // @[AxiLoadQueue.scala 163:19:@14225.4]
  wire  storeAddrNotKnownFlags_14_0; // @[AxiLoadQueue.scala 163:19:@14243.4]
  wire  storeAddrNotKnownFlags_14_1; // @[AxiLoadQueue.scala 163:19:@14245.4]
  wire  storeAddrNotKnownFlags_14_2; // @[AxiLoadQueue.scala 163:19:@14247.4]
  wire  storeAddrNotKnownFlags_14_3; // @[AxiLoadQueue.scala 163:19:@14249.4]
  wire  storeAddrNotKnownFlags_14_4; // @[AxiLoadQueue.scala 163:19:@14251.4]
  wire  storeAddrNotKnownFlags_14_5; // @[AxiLoadQueue.scala 163:19:@14253.4]
  wire  storeAddrNotKnownFlags_14_6; // @[AxiLoadQueue.scala 163:19:@14255.4]
  wire  storeAddrNotKnownFlags_14_7; // @[AxiLoadQueue.scala 163:19:@14257.4]
  wire  storeAddrNotKnownFlags_14_8; // @[AxiLoadQueue.scala 163:19:@14259.4]
  wire  storeAddrNotKnownFlags_14_9; // @[AxiLoadQueue.scala 163:19:@14261.4]
  wire  storeAddrNotKnownFlags_14_10; // @[AxiLoadQueue.scala 163:19:@14263.4]
  wire  storeAddrNotKnownFlags_14_11; // @[AxiLoadQueue.scala 163:19:@14265.4]
  wire  storeAddrNotKnownFlags_14_12; // @[AxiLoadQueue.scala 163:19:@14267.4]
  wire  storeAddrNotKnownFlags_14_13; // @[AxiLoadQueue.scala 163:19:@14269.4]
  wire  storeAddrNotKnownFlags_14_14; // @[AxiLoadQueue.scala 163:19:@14271.4]
  wire  storeAddrNotKnownFlags_14_15; // @[AxiLoadQueue.scala 163:19:@14273.4]
  wire  storeAddrNotKnownFlags_15_0; // @[AxiLoadQueue.scala 163:19:@14291.4]
  wire  storeAddrNotKnownFlags_15_1; // @[AxiLoadQueue.scala 163:19:@14293.4]
  wire  storeAddrNotKnownFlags_15_2; // @[AxiLoadQueue.scala 163:19:@14295.4]
  wire  storeAddrNotKnownFlags_15_3; // @[AxiLoadQueue.scala 163:19:@14297.4]
  wire  storeAddrNotKnownFlags_15_4; // @[AxiLoadQueue.scala 163:19:@14299.4]
  wire  storeAddrNotKnownFlags_15_5; // @[AxiLoadQueue.scala 163:19:@14301.4]
  wire  storeAddrNotKnownFlags_15_6; // @[AxiLoadQueue.scala 163:19:@14303.4]
  wire  storeAddrNotKnownFlags_15_7; // @[AxiLoadQueue.scala 163:19:@14305.4]
  wire  storeAddrNotKnownFlags_15_8; // @[AxiLoadQueue.scala 163:19:@14307.4]
  wire  storeAddrNotKnownFlags_15_9; // @[AxiLoadQueue.scala 163:19:@14309.4]
  wire  storeAddrNotKnownFlags_15_10; // @[AxiLoadQueue.scala 163:19:@14311.4]
  wire  storeAddrNotKnownFlags_15_11; // @[AxiLoadQueue.scala 163:19:@14313.4]
  wire  storeAddrNotKnownFlags_15_12; // @[AxiLoadQueue.scala 163:19:@14315.4]
  wire  storeAddrNotKnownFlags_15_13; // @[AxiLoadQueue.scala 163:19:@14317.4]
  wire  storeAddrNotKnownFlags_15_14; // @[AxiLoadQueue.scala 163:19:@14319.4]
  wire  storeAddrNotKnownFlags_15_15; // @[AxiLoadQueue.scala 163:19:@14321.4]
  wire [7:0] _T_18008; // @[Mux.scala 19:72:@14652.4]
  wire [7:0] _T_18015; // @[Mux.scala 19:72:@14659.4]
  wire [15:0] _T_18016; // @[Mux.scala 19:72:@14660.4]
  wire [15:0] _T_18018; // @[Mux.scala 19:72:@14661.4]
  wire [7:0] _T_18025; // @[Mux.scala 19:72:@14668.4]
  wire [7:0] _T_18032; // @[Mux.scala 19:72:@14675.4]
  wire [15:0] _T_18033; // @[Mux.scala 19:72:@14676.4]
  wire [15:0] _T_18035; // @[Mux.scala 19:72:@14677.4]
  wire [7:0] _T_18042; // @[Mux.scala 19:72:@14684.4]
  wire [7:0] _T_18049; // @[Mux.scala 19:72:@14691.4]
  wire [15:0] _T_18050; // @[Mux.scala 19:72:@14692.4]
  wire [15:0] _T_18052; // @[Mux.scala 19:72:@14693.4]
  wire [7:0] _T_18059; // @[Mux.scala 19:72:@14700.4]
  wire [7:0] _T_18066; // @[Mux.scala 19:72:@14707.4]
  wire [15:0] _T_18067; // @[Mux.scala 19:72:@14708.4]
  wire [15:0] _T_18069; // @[Mux.scala 19:72:@14709.4]
  wire [7:0] _T_18076; // @[Mux.scala 19:72:@14716.4]
  wire [7:0] _T_18083; // @[Mux.scala 19:72:@14723.4]
  wire [15:0] _T_18084; // @[Mux.scala 19:72:@14724.4]
  wire [15:0] _T_18086; // @[Mux.scala 19:72:@14725.4]
  wire [7:0] _T_18093; // @[Mux.scala 19:72:@14732.4]
  wire [7:0] _T_18100; // @[Mux.scala 19:72:@14739.4]
  wire [15:0] _T_18101; // @[Mux.scala 19:72:@14740.4]
  wire [15:0] _T_18103; // @[Mux.scala 19:72:@14741.4]
  wire [7:0] _T_18110; // @[Mux.scala 19:72:@14748.4]
  wire [7:0] _T_18117; // @[Mux.scala 19:72:@14755.4]
  wire [15:0] _T_18118; // @[Mux.scala 19:72:@14756.4]
  wire [15:0] _T_18120; // @[Mux.scala 19:72:@14757.4]
  wire [7:0] _T_18127; // @[Mux.scala 19:72:@14764.4]
  wire [7:0] _T_18134; // @[Mux.scala 19:72:@14771.4]
  wire [15:0] _T_18135; // @[Mux.scala 19:72:@14772.4]
  wire [15:0] _T_18137; // @[Mux.scala 19:72:@14773.4]
  wire [15:0] _T_18152; // @[Mux.scala 19:72:@14788.4]
  wire [15:0] _T_18154; // @[Mux.scala 19:72:@14789.4]
  wire [15:0] _T_18169; // @[Mux.scala 19:72:@14804.4]
  wire [15:0] _T_18171; // @[Mux.scala 19:72:@14805.4]
  wire [15:0] _T_18186; // @[Mux.scala 19:72:@14820.4]
  wire [15:0] _T_18188; // @[Mux.scala 19:72:@14821.4]
  wire [15:0] _T_18203; // @[Mux.scala 19:72:@14836.4]
  wire [15:0] _T_18205; // @[Mux.scala 19:72:@14837.4]
  wire [15:0] _T_18220; // @[Mux.scala 19:72:@14852.4]
  wire [15:0] _T_18222; // @[Mux.scala 19:72:@14853.4]
  wire [15:0] _T_18237; // @[Mux.scala 19:72:@14868.4]
  wire [15:0] _T_18239; // @[Mux.scala 19:72:@14869.4]
  wire [15:0] _T_18254; // @[Mux.scala 19:72:@14884.4]
  wire [15:0] _T_18256; // @[Mux.scala 19:72:@14885.4]
  wire [15:0] _T_18271; // @[Mux.scala 19:72:@14900.4]
  wire [15:0] _T_18273; // @[Mux.scala 19:72:@14901.4]
  wire [15:0] _T_18274; // @[Mux.scala 19:72:@14902.4]
  wire [15:0] _T_18275; // @[Mux.scala 19:72:@14903.4]
  wire [15:0] _T_18276; // @[Mux.scala 19:72:@14904.4]
  wire [15:0] _T_18277; // @[Mux.scala 19:72:@14905.4]
  wire [15:0] _T_18278; // @[Mux.scala 19:72:@14906.4]
  wire [15:0] _T_18279; // @[Mux.scala 19:72:@14907.4]
  wire [15:0] _T_18280; // @[Mux.scala 19:72:@14908.4]
  wire [15:0] _T_18281; // @[Mux.scala 19:72:@14909.4]
  wire [15:0] _T_18282; // @[Mux.scala 19:72:@14910.4]
  wire [15:0] _T_18283; // @[Mux.scala 19:72:@14911.4]
  wire [15:0] _T_18284; // @[Mux.scala 19:72:@14912.4]
  wire [15:0] _T_18285; // @[Mux.scala 19:72:@14913.4]
  wire [15:0] _T_18286; // @[Mux.scala 19:72:@14914.4]
  wire [15:0] _T_18287; // @[Mux.scala 19:72:@14915.4]
  wire [15:0] _T_18288; // @[Mux.scala 19:72:@14916.4]
  wire [7:0] _T_18866; // @[Mux.scala 19:72:@15266.4]
  wire [7:0] _T_18873; // @[Mux.scala 19:72:@15273.4]
  wire [15:0] _T_18874; // @[Mux.scala 19:72:@15274.4]
  wire [15:0] _T_18876; // @[Mux.scala 19:72:@15275.4]
  wire [7:0] _T_18883; // @[Mux.scala 19:72:@15282.4]
  wire [7:0] _T_18890; // @[Mux.scala 19:72:@15289.4]
  wire [15:0] _T_18891; // @[Mux.scala 19:72:@15290.4]
  wire [15:0] _T_18893; // @[Mux.scala 19:72:@15291.4]
  wire [7:0] _T_18900; // @[Mux.scala 19:72:@15298.4]
  wire [7:0] _T_18907; // @[Mux.scala 19:72:@15305.4]
  wire [15:0] _T_18908; // @[Mux.scala 19:72:@15306.4]
  wire [15:0] _T_18910; // @[Mux.scala 19:72:@15307.4]
  wire [7:0] _T_18917; // @[Mux.scala 19:72:@15314.4]
  wire [7:0] _T_18924; // @[Mux.scala 19:72:@15321.4]
  wire [15:0] _T_18925; // @[Mux.scala 19:72:@15322.4]
  wire [15:0] _T_18927; // @[Mux.scala 19:72:@15323.4]
  wire [7:0] _T_18934; // @[Mux.scala 19:72:@15330.4]
  wire [7:0] _T_18941; // @[Mux.scala 19:72:@15337.4]
  wire [15:0] _T_18942; // @[Mux.scala 19:72:@15338.4]
  wire [15:0] _T_18944; // @[Mux.scala 19:72:@15339.4]
  wire [7:0] _T_18951; // @[Mux.scala 19:72:@15346.4]
  wire [7:0] _T_18958; // @[Mux.scala 19:72:@15353.4]
  wire [15:0] _T_18959; // @[Mux.scala 19:72:@15354.4]
  wire [15:0] _T_18961; // @[Mux.scala 19:72:@15355.4]
  wire [7:0] _T_18968; // @[Mux.scala 19:72:@15362.4]
  wire [7:0] _T_18975; // @[Mux.scala 19:72:@15369.4]
  wire [15:0] _T_18976; // @[Mux.scala 19:72:@15370.4]
  wire [15:0] _T_18978; // @[Mux.scala 19:72:@15371.4]
  wire [7:0] _T_18985; // @[Mux.scala 19:72:@15378.4]
  wire [7:0] _T_18992; // @[Mux.scala 19:72:@15385.4]
  wire [15:0] _T_18993; // @[Mux.scala 19:72:@15386.4]
  wire [15:0] _T_18995; // @[Mux.scala 19:72:@15387.4]
  wire [15:0] _T_19010; // @[Mux.scala 19:72:@15402.4]
  wire [15:0] _T_19012; // @[Mux.scala 19:72:@15403.4]
  wire [15:0] _T_19027; // @[Mux.scala 19:72:@15418.4]
  wire [15:0] _T_19029; // @[Mux.scala 19:72:@15419.4]
  wire [15:0] _T_19044; // @[Mux.scala 19:72:@15434.4]
  wire [15:0] _T_19046; // @[Mux.scala 19:72:@15435.4]
  wire [15:0] _T_19061; // @[Mux.scala 19:72:@15450.4]
  wire [15:0] _T_19063; // @[Mux.scala 19:72:@15451.4]
  wire [15:0] _T_19078; // @[Mux.scala 19:72:@15466.4]
  wire [15:0] _T_19080; // @[Mux.scala 19:72:@15467.4]
  wire [15:0] _T_19095; // @[Mux.scala 19:72:@15482.4]
  wire [15:0] _T_19097; // @[Mux.scala 19:72:@15483.4]
  wire [15:0] _T_19112; // @[Mux.scala 19:72:@15498.4]
  wire [15:0] _T_19114; // @[Mux.scala 19:72:@15499.4]
  wire [15:0] _T_19129; // @[Mux.scala 19:72:@15514.4]
  wire [15:0] _T_19131; // @[Mux.scala 19:72:@15515.4]
  wire [15:0] _T_19132; // @[Mux.scala 19:72:@15516.4]
  wire [15:0] _T_19133; // @[Mux.scala 19:72:@15517.4]
  wire [15:0] _T_19134; // @[Mux.scala 19:72:@15518.4]
  wire [15:0] _T_19135; // @[Mux.scala 19:72:@15519.4]
  wire [15:0] _T_19136; // @[Mux.scala 19:72:@15520.4]
  wire [15:0] _T_19137; // @[Mux.scala 19:72:@15521.4]
  wire [15:0] _T_19138; // @[Mux.scala 19:72:@15522.4]
  wire [15:0] _T_19139; // @[Mux.scala 19:72:@15523.4]
  wire [15:0] _T_19140; // @[Mux.scala 19:72:@15524.4]
  wire [15:0] _T_19141; // @[Mux.scala 19:72:@15525.4]
  wire [15:0] _T_19142; // @[Mux.scala 19:72:@15526.4]
  wire [15:0] _T_19143; // @[Mux.scala 19:72:@15527.4]
  wire [15:0] _T_19144; // @[Mux.scala 19:72:@15528.4]
  wire [15:0] _T_19145; // @[Mux.scala 19:72:@15529.4]
  wire [15:0] _T_19146; // @[Mux.scala 19:72:@15530.4]
  wire [7:0] _T_19724; // @[Mux.scala 19:72:@15880.4]
  wire [7:0] _T_19731; // @[Mux.scala 19:72:@15887.4]
  wire [15:0] _T_19732; // @[Mux.scala 19:72:@15888.4]
  wire [15:0] _T_19734; // @[Mux.scala 19:72:@15889.4]
  wire [7:0] _T_19741; // @[Mux.scala 19:72:@15896.4]
  wire [7:0] _T_19748; // @[Mux.scala 19:72:@15903.4]
  wire [15:0] _T_19749; // @[Mux.scala 19:72:@15904.4]
  wire [15:0] _T_19751; // @[Mux.scala 19:72:@15905.4]
  wire [7:0] _T_19758; // @[Mux.scala 19:72:@15912.4]
  wire [7:0] _T_19765; // @[Mux.scala 19:72:@15919.4]
  wire [15:0] _T_19766; // @[Mux.scala 19:72:@15920.4]
  wire [15:0] _T_19768; // @[Mux.scala 19:72:@15921.4]
  wire [7:0] _T_19775; // @[Mux.scala 19:72:@15928.4]
  wire [7:0] _T_19782; // @[Mux.scala 19:72:@15935.4]
  wire [15:0] _T_19783; // @[Mux.scala 19:72:@15936.4]
  wire [15:0] _T_19785; // @[Mux.scala 19:72:@15937.4]
  wire [7:0] _T_19792; // @[Mux.scala 19:72:@15944.4]
  wire [7:0] _T_19799; // @[Mux.scala 19:72:@15951.4]
  wire [15:0] _T_19800; // @[Mux.scala 19:72:@15952.4]
  wire [15:0] _T_19802; // @[Mux.scala 19:72:@15953.4]
  wire [7:0] _T_19809; // @[Mux.scala 19:72:@15960.4]
  wire [7:0] _T_19816; // @[Mux.scala 19:72:@15967.4]
  wire [15:0] _T_19817; // @[Mux.scala 19:72:@15968.4]
  wire [15:0] _T_19819; // @[Mux.scala 19:72:@15969.4]
  wire [7:0] _T_19826; // @[Mux.scala 19:72:@15976.4]
  wire [7:0] _T_19833; // @[Mux.scala 19:72:@15983.4]
  wire [15:0] _T_19834; // @[Mux.scala 19:72:@15984.4]
  wire [15:0] _T_19836; // @[Mux.scala 19:72:@15985.4]
  wire [7:0] _T_19843; // @[Mux.scala 19:72:@15992.4]
  wire [7:0] _T_19850; // @[Mux.scala 19:72:@15999.4]
  wire [15:0] _T_19851; // @[Mux.scala 19:72:@16000.4]
  wire [15:0] _T_19853; // @[Mux.scala 19:72:@16001.4]
  wire [15:0] _T_19868; // @[Mux.scala 19:72:@16016.4]
  wire [15:0] _T_19870; // @[Mux.scala 19:72:@16017.4]
  wire [15:0] _T_19885; // @[Mux.scala 19:72:@16032.4]
  wire [15:0] _T_19887; // @[Mux.scala 19:72:@16033.4]
  wire [15:0] _T_19902; // @[Mux.scala 19:72:@16048.4]
  wire [15:0] _T_19904; // @[Mux.scala 19:72:@16049.4]
  wire [15:0] _T_19919; // @[Mux.scala 19:72:@16064.4]
  wire [15:0] _T_19921; // @[Mux.scala 19:72:@16065.4]
  wire [15:0] _T_19936; // @[Mux.scala 19:72:@16080.4]
  wire [15:0] _T_19938; // @[Mux.scala 19:72:@16081.4]
  wire [15:0] _T_19953; // @[Mux.scala 19:72:@16096.4]
  wire [15:0] _T_19955; // @[Mux.scala 19:72:@16097.4]
  wire [15:0] _T_19970; // @[Mux.scala 19:72:@16112.4]
  wire [15:0] _T_19972; // @[Mux.scala 19:72:@16113.4]
  wire [15:0] _T_19987; // @[Mux.scala 19:72:@16128.4]
  wire [15:0] _T_19989; // @[Mux.scala 19:72:@16129.4]
  wire [15:0] _T_19990; // @[Mux.scala 19:72:@16130.4]
  wire [15:0] _T_19991; // @[Mux.scala 19:72:@16131.4]
  wire [15:0] _T_19992; // @[Mux.scala 19:72:@16132.4]
  wire [15:0] _T_19993; // @[Mux.scala 19:72:@16133.4]
  wire [15:0] _T_19994; // @[Mux.scala 19:72:@16134.4]
  wire [15:0] _T_19995; // @[Mux.scala 19:72:@16135.4]
  wire [15:0] _T_19996; // @[Mux.scala 19:72:@16136.4]
  wire [15:0] _T_19997; // @[Mux.scala 19:72:@16137.4]
  wire [15:0] _T_19998; // @[Mux.scala 19:72:@16138.4]
  wire [15:0] _T_19999; // @[Mux.scala 19:72:@16139.4]
  wire [15:0] _T_20000; // @[Mux.scala 19:72:@16140.4]
  wire [15:0] _T_20001; // @[Mux.scala 19:72:@16141.4]
  wire [15:0] _T_20002; // @[Mux.scala 19:72:@16142.4]
  wire [15:0] _T_20003; // @[Mux.scala 19:72:@16143.4]
  wire [15:0] _T_20004; // @[Mux.scala 19:72:@16144.4]
  wire [7:0] _T_20582; // @[Mux.scala 19:72:@16494.4]
  wire [7:0] _T_20589; // @[Mux.scala 19:72:@16501.4]
  wire [15:0] _T_20590; // @[Mux.scala 19:72:@16502.4]
  wire [15:0] _T_20592; // @[Mux.scala 19:72:@16503.4]
  wire [7:0] _T_20599; // @[Mux.scala 19:72:@16510.4]
  wire [7:0] _T_20606; // @[Mux.scala 19:72:@16517.4]
  wire [15:0] _T_20607; // @[Mux.scala 19:72:@16518.4]
  wire [15:0] _T_20609; // @[Mux.scala 19:72:@16519.4]
  wire [7:0] _T_20616; // @[Mux.scala 19:72:@16526.4]
  wire [7:0] _T_20623; // @[Mux.scala 19:72:@16533.4]
  wire [15:0] _T_20624; // @[Mux.scala 19:72:@16534.4]
  wire [15:0] _T_20626; // @[Mux.scala 19:72:@16535.4]
  wire [7:0] _T_20633; // @[Mux.scala 19:72:@16542.4]
  wire [7:0] _T_20640; // @[Mux.scala 19:72:@16549.4]
  wire [15:0] _T_20641; // @[Mux.scala 19:72:@16550.4]
  wire [15:0] _T_20643; // @[Mux.scala 19:72:@16551.4]
  wire [7:0] _T_20650; // @[Mux.scala 19:72:@16558.4]
  wire [7:0] _T_20657; // @[Mux.scala 19:72:@16565.4]
  wire [15:0] _T_20658; // @[Mux.scala 19:72:@16566.4]
  wire [15:0] _T_20660; // @[Mux.scala 19:72:@16567.4]
  wire [7:0] _T_20667; // @[Mux.scala 19:72:@16574.4]
  wire [7:0] _T_20674; // @[Mux.scala 19:72:@16581.4]
  wire [15:0] _T_20675; // @[Mux.scala 19:72:@16582.4]
  wire [15:0] _T_20677; // @[Mux.scala 19:72:@16583.4]
  wire [7:0] _T_20684; // @[Mux.scala 19:72:@16590.4]
  wire [7:0] _T_20691; // @[Mux.scala 19:72:@16597.4]
  wire [15:0] _T_20692; // @[Mux.scala 19:72:@16598.4]
  wire [15:0] _T_20694; // @[Mux.scala 19:72:@16599.4]
  wire [7:0] _T_20701; // @[Mux.scala 19:72:@16606.4]
  wire [7:0] _T_20708; // @[Mux.scala 19:72:@16613.4]
  wire [15:0] _T_20709; // @[Mux.scala 19:72:@16614.4]
  wire [15:0] _T_20711; // @[Mux.scala 19:72:@16615.4]
  wire [15:0] _T_20726; // @[Mux.scala 19:72:@16630.4]
  wire [15:0] _T_20728; // @[Mux.scala 19:72:@16631.4]
  wire [15:0] _T_20743; // @[Mux.scala 19:72:@16646.4]
  wire [15:0] _T_20745; // @[Mux.scala 19:72:@16647.4]
  wire [15:0] _T_20760; // @[Mux.scala 19:72:@16662.4]
  wire [15:0] _T_20762; // @[Mux.scala 19:72:@16663.4]
  wire [15:0] _T_20777; // @[Mux.scala 19:72:@16678.4]
  wire [15:0] _T_20779; // @[Mux.scala 19:72:@16679.4]
  wire [15:0] _T_20794; // @[Mux.scala 19:72:@16694.4]
  wire [15:0] _T_20796; // @[Mux.scala 19:72:@16695.4]
  wire [15:0] _T_20811; // @[Mux.scala 19:72:@16710.4]
  wire [15:0] _T_20813; // @[Mux.scala 19:72:@16711.4]
  wire [15:0] _T_20828; // @[Mux.scala 19:72:@16726.4]
  wire [15:0] _T_20830; // @[Mux.scala 19:72:@16727.4]
  wire [15:0] _T_20845; // @[Mux.scala 19:72:@16742.4]
  wire [15:0] _T_20847; // @[Mux.scala 19:72:@16743.4]
  wire [15:0] _T_20848; // @[Mux.scala 19:72:@16744.4]
  wire [15:0] _T_20849; // @[Mux.scala 19:72:@16745.4]
  wire [15:0] _T_20850; // @[Mux.scala 19:72:@16746.4]
  wire [15:0] _T_20851; // @[Mux.scala 19:72:@16747.4]
  wire [15:0] _T_20852; // @[Mux.scala 19:72:@16748.4]
  wire [15:0] _T_20853; // @[Mux.scala 19:72:@16749.4]
  wire [15:0] _T_20854; // @[Mux.scala 19:72:@16750.4]
  wire [15:0] _T_20855; // @[Mux.scala 19:72:@16751.4]
  wire [15:0] _T_20856; // @[Mux.scala 19:72:@16752.4]
  wire [15:0] _T_20857; // @[Mux.scala 19:72:@16753.4]
  wire [15:0] _T_20858; // @[Mux.scala 19:72:@16754.4]
  wire [15:0] _T_20859; // @[Mux.scala 19:72:@16755.4]
  wire [15:0] _T_20860; // @[Mux.scala 19:72:@16756.4]
  wire [15:0] _T_20861; // @[Mux.scala 19:72:@16757.4]
  wire [15:0] _T_20862; // @[Mux.scala 19:72:@16758.4]
  wire [7:0] _T_21440; // @[Mux.scala 19:72:@17108.4]
  wire [7:0] _T_21447; // @[Mux.scala 19:72:@17115.4]
  wire [15:0] _T_21448; // @[Mux.scala 19:72:@17116.4]
  wire [15:0] _T_21450; // @[Mux.scala 19:72:@17117.4]
  wire [7:0] _T_21457; // @[Mux.scala 19:72:@17124.4]
  wire [7:0] _T_21464; // @[Mux.scala 19:72:@17131.4]
  wire [15:0] _T_21465; // @[Mux.scala 19:72:@17132.4]
  wire [15:0] _T_21467; // @[Mux.scala 19:72:@17133.4]
  wire [7:0] _T_21474; // @[Mux.scala 19:72:@17140.4]
  wire [7:0] _T_21481; // @[Mux.scala 19:72:@17147.4]
  wire [15:0] _T_21482; // @[Mux.scala 19:72:@17148.4]
  wire [15:0] _T_21484; // @[Mux.scala 19:72:@17149.4]
  wire [7:0] _T_21491; // @[Mux.scala 19:72:@17156.4]
  wire [7:0] _T_21498; // @[Mux.scala 19:72:@17163.4]
  wire [15:0] _T_21499; // @[Mux.scala 19:72:@17164.4]
  wire [15:0] _T_21501; // @[Mux.scala 19:72:@17165.4]
  wire [7:0] _T_21508; // @[Mux.scala 19:72:@17172.4]
  wire [7:0] _T_21515; // @[Mux.scala 19:72:@17179.4]
  wire [15:0] _T_21516; // @[Mux.scala 19:72:@17180.4]
  wire [15:0] _T_21518; // @[Mux.scala 19:72:@17181.4]
  wire [7:0] _T_21525; // @[Mux.scala 19:72:@17188.4]
  wire [7:0] _T_21532; // @[Mux.scala 19:72:@17195.4]
  wire [15:0] _T_21533; // @[Mux.scala 19:72:@17196.4]
  wire [15:0] _T_21535; // @[Mux.scala 19:72:@17197.4]
  wire [7:0] _T_21542; // @[Mux.scala 19:72:@17204.4]
  wire [7:0] _T_21549; // @[Mux.scala 19:72:@17211.4]
  wire [15:0] _T_21550; // @[Mux.scala 19:72:@17212.4]
  wire [15:0] _T_21552; // @[Mux.scala 19:72:@17213.4]
  wire [7:0] _T_21559; // @[Mux.scala 19:72:@17220.4]
  wire [7:0] _T_21566; // @[Mux.scala 19:72:@17227.4]
  wire [15:0] _T_21567; // @[Mux.scala 19:72:@17228.4]
  wire [15:0] _T_21569; // @[Mux.scala 19:72:@17229.4]
  wire [15:0] _T_21584; // @[Mux.scala 19:72:@17244.4]
  wire [15:0] _T_21586; // @[Mux.scala 19:72:@17245.4]
  wire [15:0] _T_21601; // @[Mux.scala 19:72:@17260.4]
  wire [15:0] _T_21603; // @[Mux.scala 19:72:@17261.4]
  wire [15:0] _T_21618; // @[Mux.scala 19:72:@17276.4]
  wire [15:0] _T_21620; // @[Mux.scala 19:72:@17277.4]
  wire [15:0] _T_21635; // @[Mux.scala 19:72:@17292.4]
  wire [15:0] _T_21637; // @[Mux.scala 19:72:@17293.4]
  wire [15:0] _T_21652; // @[Mux.scala 19:72:@17308.4]
  wire [15:0] _T_21654; // @[Mux.scala 19:72:@17309.4]
  wire [15:0] _T_21669; // @[Mux.scala 19:72:@17324.4]
  wire [15:0] _T_21671; // @[Mux.scala 19:72:@17325.4]
  wire [15:0] _T_21686; // @[Mux.scala 19:72:@17340.4]
  wire [15:0] _T_21688; // @[Mux.scala 19:72:@17341.4]
  wire [15:0] _T_21703; // @[Mux.scala 19:72:@17356.4]
  wire [15:0] _T_21705; // @[Mux.scala 19:72:@17357.4]
  wire [15:0] _T_21706; // @[Mux.scala 19:72:@17358.4]
  wire [15:0] _T_21707; // @[Mux.scala 19:72:@17359.4]
  wire [15:0] _T_21708; // @[Mux.scala 19:72:@17360.4]
  wire [15:0] _T_21709; // @[Mux.scala 19:72:@17361.4]
  wire [15:0] _T_21710; // @[Mux.scala 19:72:@17362.4]
  wire [15:0] _T_21711; // @[Mux.scala 19:72:@17363.4]
  wire [15:0] _T_21712; // @[Mux.scala 19:72:@17364.4]
  wire [15:0] _T_21713; // @[Mux.scala 19:72:@17365.4]
  wire [15:0] _T_21714; // @[Mux.scala 19:72:@17366.4]
  wire [15:0] _T_21715; // @[Mux.scala 19:72:@17367.4]
  wire [15:0] _T_21716; // @[Mux.scala 19:72:@17368.4]
  wire [15:0] _T_21717; // @[Mux.scala 19:72:@17369.4]
  wire [15:0] _T_21718; // @[Mux.scala 19:72:@17370.4]
  wire [15:0] _T_21719; // @[Mux.scala 19:72:@17371.4]
  wire [15:0] _T_21720; // @[Mux.scala 19:72:@17372.4]
  wire [7:0] _T_22298; // @[Mux.scala 19:72:@17722.4]
  wire [7:0] _T_22305; // @[Mux.scala 19:72:@17729.4]
  wire [15:0] _T_22306; // @[Mux.scala 19:72:@17730.4]
  wire [15:0] _T_22308; // @[Mux.scala 19:72:@17731.4]
  wire [7:0] _T_22315; // @[Mux.scala 19:72:@17738.4]
  wire [7:0] _T_22322; // @[Mux.scala 19:72:@17745.4]
  wire [15:0] _T_22323; // @[Mux.scala 19:72:@17746.4]
  wire [15:0] _T_22325; // @[Mux.scala 19:72:@17747.4]
  wire [7:0] _T_22332; // @[Mux.scala 19:72:@17754.4]
  wire [7:0] _T_22339; // @[Mux.scala 19:72:@17761.4]
  wire [15:0] _T_22340; // @[Mux.scala 19:72:@17762.4]
  wire [15:0] _T_22342; // @[Mux.scala 19:72:@17763.4]
  wire [7:0] _T_22349; // @[Mux.scala 19:72:@17770.4]
  wire [7:0] _T_22356; // @[Mux.scala 19:72:@17777.4]
  wire [15:0] _T_22357; // @[Mux.scala 19:72:@17778.4]
  wire [15:0] _T_22359; // @[Mux.scala 19:72:@17779.4]
  wire [7:0] _T_22366; // @[Mux.scala 19:72:@17786.4]
  wire [7:0] _T_22373; // @[Mux.scala 19:72:@17793.4]
  wire [15:0] _T_22374; // @[Mux.scala 19:72:@17794.4]
  wire [15:0] _T_22376; // @[Mux.scala 19:72:@17795.4]
  wire [7:0] _T_22383; // @[Mux.scala 19:72:@17802.4]
  wire [7:0] _T_22390; // @[Mux.scala 19:72:@17809.4]
  wire [15:0] _T_22391; // @[Mux.scala 19:72:@17810.4]
  wire [15:0] _T_22393; // @[Mux.scala 19:72:@17811.4]
  wire [7:0] _T_22400; // @[Mux.scala 19:72:@17818.4]
  wire [7:0] _T_22407; // @[Mux.scala 19:72:@17825.4]
  wire [15:0] _T_22408; // @[Mux.scala 19:72:@17826.4]
  wire [15:0] _T_22410; // @[Mux.scala 19:72:@17827.4]
  wire [7:0] _T_22417; // @[Mux.scala 19:72:@17834.4]
  wire [7:0] _T_22424; // @[Mux.scala 19:72:@17841.4]
  wire [15:0] _T_22425; // @[Mux.scala 19:72:@17842.4]
  wire [15:0] _T_22427; // @[Mux.scala 19:72:@17843.4]
  wire [15:0] _T_22442; // @[Mux.scala 19:72:@17858.4]
  wire [15:0] _T_22444; // @[Mux.scala 19:72:@17859.4]
  wire [15:0] _T_22459; // @[Mux.scala 19:72:@17874.4]
  wire [15:0] _T_22461; // @[Mux.scala 19:72:@17875.4]
  wire [15:0] _T_22476; // @[Mux.scala 19:72:@17890.4]
  wire [15:0] _T_22478; // @[Mux.scala 19:72:@17891.4]
  wire [15:0] _T_22493; // @[Mux.scala 19:72:@17906.4]
  wire [15:0] _T_22495; // @[Mux.scala 19:72:@17907.4]
  wire [15:0] _T_22510; // @[Mux.scala 19:72:@17922.4]
  wire [15:0] _T_22512; // @[Mux.scala 19:72:@17923.4]
  wire [15:0] _T_22527; // @[Mux.scala 19:72:@17938.4]
  wire [15:0] _T_22529; // @[Mux.scala 19:72:@17939.4]
  wire [15:0] _T_22544; // @[Mux.scala 19:72:@17954.4]
  wire [15:0] _T_22546; // @[Mux.scala 19:72:@17955.4]
  wire [15:0] _T_22561; // @[Mux.scala 19:72:@17970.4]
  wire [15:0] _T_22563; // @[Mux.scala 19:72:@17971.4]
  wire [15:0] _T_22564; // @[Mux.scala 19:72:@17972.4]
  wire [15:0] _T_22565; // @[Mux.scala 19:72:@17973.4]
  wire [15:0] _T_22566; // @[Mux.scala 19:72:@17974.4]
  wire [15:0] _T_22567; // @[Mux.scala 19:72:@17975.4]
  wire [15:0] _T_22568; // @[Mux.scala 19:72:@17976.4]
  wire [15:0] _T_22569; // @[Mux.scala 19:72:@17977.4]
  wire [15:0] _T_22570; // @[Mux.scala 19:72:@17978.4]
  wire [15:0] _T_22571; // @[Mux.scala 19:72:@17979.4]
  wire [15:0] _T_22572; // @[Mux.scala 19:72:@17980.4]
  wire [15:0] _T_22573; // @[Mux.scala 19:72:@17981.4]
  wire [15:0] _T_22574; // @[Mux.scala 19:72:@17982.4]
  wire [15:0] _T_22575; // @[Mux.scala 19:72:@17983.4]
  wire [15:0] _T_22576; // @[Mux.scala 19:72:@17984.4]
  wire [15:0] _T_22577; // @[Mux.scala 19:72:@17985.4]
  wire [15:0] _T_22578; // @[Mux.scala 19:72:@17986.4]
  wire [7:0] _T_23156; // @[Mux.scala 19:72:@18336.4]
  wire [7:0] _T_23163; // @[Mux.scala 19:72:@18343.4]
  wire [15:0] _T_23164; // @[Mux.scala 19:72:@18344.4]
  wire [15:0] _T_23166; // @[Mux.scala 19:72:@18345.4]
  wire [7:0] _T_23173; // @[Mux.scala 19:72:@18352.4]
  wire [7:0] _T_23180; // @[Mux.scala 19:72:@18359.4]
  wire [15:0] _T_23181; // @[Mux.scala 19:72:@18360.4]
  wire [15:0] _T_23183; // @[Mux.scala 19:72:@18361.4]
  wire [7:0] _T_23190; // @[Mux.scala 19:72:@18368.4]
  wire [7:0] _T_23197; // @[Mux.scala 19:72:@18375.4]
  wire [15:0] _T_23198; // @[Mux.scala 19:72:@18376.4]
  wire [15:0] _T_23200; // @[Mux.scala 19:72:@18377.4]
  wire [7:0] _T_23207; // @[Mux.scala 19:72:@18384.4]
  wire [7:0] _T_23214; // @[Mux.scala 19:72:@18391.4]
  wire [15:0] _T_23215; // @[Mux.scala 19:72:@18392.4]
  wire [15:0] _T_23217; // @[Mux.scala 19:72:@18393.4]
  wire [7:0] _T_23224; // @[Mux.scala 19:72:@18400.4]
  wire [7:0] _T_23231; // @[Mux.scala 19:72:@18407.4]
  wire [15:0] _T_23232; // @[Mux.scala 19:72:@18408.4]
  wire [15:0] _T_23234; // @[Mux.scala 19:72:@18409.4]
  wire [7:0] _T_23241; // @[Mux.scala 19:72:@18416.4]
  wire [7:0] _T_23248; // @[Mux.scala 19:72:@18423.4]
  wire [15:0] _T_23249; // @[Mux.scala 19:72:@18424.4]
  wire [15:0] _T_23251; // @[Mux.scala 19:72:@18425.4]
  wire [7:0] _T_23258; // @[Mux.scala 19:72:@18432.4]
  wire [7:0] _T_23265; // @[Mux.scala 19:72:@18439.4]
  wire [15:0] _T_23266; // @[Mux.scala 19:72:@18440.4]
  wire [15:0] _T_23268; // @[Mux.scala 19:72:@18441.4]
  wire [7:0] _T_23275; // @[Mux.scala 19:72:@18448.4]
  wire [7:0] _T_23282; // @[Mux.scala 19:72:@18455.4]
  wire [15:0] _T_23283; // @[Mux.scala 19:72:@18456.4]
  wire [15:0] _T_23285; // @[Mux.scala 19:72:@18457.4]
  wire [15:0] _T_23300; // @[Mux.scala 19:72:@18472.4]
  wire [15:0] _T_23302; // @[Mux.scala 19:72:@18473.4]
  wire [15:0] _T_23317; // @[Mux.scala 19:72:@18488.4]
  wire [15:0] _T_23319; // @[Mux.scala 19:72:@18489.4]
  wire [15:0] _T_23334; // @[Mux.scala 19:72:@18504.4]
  wire [15:0] _T_23336; // @[Mux.scala 19:72:@18505.4]
  wire [15:0] _T_23351; // @[Mux.scala 19:72:@18520.4]
  wire [15:0] _T_23353; // @[Mux.scala 19:72:@18521.4]
  wire [15:0] _T_23368; // @[Mux.scala 19:72:@18536.4]
  wire [15:0] _T_23370; // @[Mux.scala 19:72:@18537.4]
  wire [15:0] _T_23385; // @[Mux.scala 19:72:@18552.4]
  wire [15:0] _T_23387; // @[Mux.scala 19:72:@18553.4]
  wire [15:0] _T_23402; // @[Mux.scala 19:72:@18568.4]
  wire [15:0] _T_23404; // @[Mux.scala 19:72:@18569.4]
  wire [15:0] _T_23419; // @[Mux.scala 19:72:@18584.4]
  wire [15:0] _T_23421; // @[Mux.scala 19:72:@18585.4]
  wire [15:0] _T_23422; // @[Mux.scala 19:72:@18586.4]
  wire [15:0] _T_23423; // @[Mux.scala 19:72:@18587.4]
  wire [15:0] _T_23424; // @[Mux.scala 19:72:@18588.4]
  wire [15:0] _T_23425; // @[Mux.scala 19:72:@18589.4]
  wire [15:0] _T_23426; // @[Mux.scala 19:72:@18590.4]
  wire [15:0] _T_23427; // @[Mux.scala 19:72:@18591.4]
  wire [15:0] _T_23428; // @[Mux.scala 19:72:@18592.4]
  wire [15:0] _T_23429; // @[Mux.scala 19:72:@18593.4]
  wire [15:0] _T_23430; // @[Mux.scala 19:72:@18594.4]
  wire [15:0] _T_23431; // @[Mux.scala 19:72:@18595.4]
  wire [15:0] _T_23432; // @[Mux.scala 19:72:@18596.4]
  wire [15:0] _T_23433; // @[Mux.scala 19:72:@18597.4]
  wire [15:0] _T_23434; // @[Mux.scala 19:72:@18598.4]
  wire [15:0] _T_23435; // @[Mux.scala 19:72:@18599.4]
  wire [15:0] _T_23436; // @[Mux.scala 19:72:@18600.4]
  wire [7:0] _T_24014; // @[Mux.scala 19:72:@18950.4]
  wire [7:0] _T_24021; // @[Mux.scala 19:72:@18957.4]
  wire [15:0] _T_24022; // @[Mux.scala 19:72:@18958.4]
  wire [15:0] _T_24024; // @[Mux.scala 19:72:@18959.4]
  wire [7:0] _T_24031; // @[Mux.scala 19:72:@18966.4]
  wire [7:0] _T_24038; // @[Mux.scala 19:72:@18973.4]
  wire [15:0] _T_24039; // @[Mux.scala 19:72:@18974.4]
  wire [15:0] _T_24041; // @[Mux.scala 19:72:@18975.4]
  wire [7:0] _T_24048; // @[Mux.scala 19:72:@18982.4]
  wire [7:0] _T_24055; // @[Mux.scala 19:72:@18989.4]
  wire [15:0] _T_24056; // @[Mux.scala 19:72:@18990.4]
  wire [15:0] _T_24058; // @[Mux.scala 19:72:@18991.4]
  wire [7:0] _T_24065; // @[Mux.scala 19:72:@18998.4]
  wire [7:0] _T_24072; // @[Mux.scala 19:72:@19005.4]
  wire [15:0] _T_24073; // @[Mux.scala 19:72:@19006.4]
  wire [15:0] _T_24075; // @[Mux.scala 19:72:@19007.4]
  wire [7:0] _T_24082; // @[Mux.scala 19:72:@19014.4]
  wire [7:0] _T_24089; // @[Mux.scala 19:72:@19021.4]
  wire [15:0] _T_24090; // @[Mux.scala 19:72:@19022.4]
  wire [15:0] _T_24092; // @[Mux.scala 19:72:@19023.4]
  wire [7:0] _T_24099; // @[Mux.scala 19:72:@19030.4]
  wire [7:0] _T_24106; // @[Mux.scala 19:72:@19037.4]
  wire [15:0] _T_24107; // @[Mux.scala 19:72:@19038.4]
  wire [15:0] _T_24109; // @[Mux.scala 19:72:@19039.4]
  wire [7:0] _T_24116; // @[Mux.scala 19:72:@19046.4]
  wire [7:0] _T_24123; // @[Mux.scala 19:72:@19053.4]
  wire [15:0] _T_24124; // @[Mux.scala 19:72:@19054.4]
  wire [15:0] _T_24126; // @[Mux.scala 19:72:@19055.4]
  wire [7:0] _T_24133; // @[Mux.scala 19:72:@19062.4]
  wire [7:0] _T_24140; // @[Mux.scala 19:72:@19069.4]
  wire [15:0] _T_24141; // @[Mux.scala 19:72:@19070.4]
  wire [15:0] _T_24143; // @[Mux.scala 19:72:@19071.4]
  wire [15:0] _T_24158; // @[Mux.scala 19:72:@19086.4]
  wire [15:0] _T_24160; // @[Mux.scala 19:72:@19087.4]
  wire [15:0] _T_24175; // @[Mux.scala 19:72:@19102.4]
  wire [15:0] _T_24177; // @[Mux.scala 19:72:@19103.4]
  wire [15:0] _T_24192; // @[Mux.scala 19:72:@19118.4]
  wire [15:0] _T_24194; // @[Mux.scala 19:72:@19119.4]
  wire [15:0] _T_24209; // @[Mux.scala 19:72:@19134.4]
  wire [15:0] _T_24211; // @[Mux.scala 19:72:@19135.4]
  wire [15:0] _T_24226; // @[Mux.scala 19:72:@19150.4]
  wire [15:0] _T_24228; // @[Mux.scala 19:72:@19151.4]
  wire [15:0] _T_24243; // @[Mux.scala 19:72:@19166.4]
  wire [15:0] _T_24245; // @[Mux.scala 19:72:@19167.4]
  wire [15:0] _T_24260; // @[Mux.scala 19:72:@19182.4]
  wire [15:0] _T_24262; // @[Mux.scala 19:72:@19183.4]
  wire [15:0] _T_24277; // @[Mux.scala 19:72:@19198.4]
  wire [15:0] _T_24279; // @[Mux.scala 19:72:@19199.4]
  wire [15:0] _T_24280; // @[Mux.scala 19:72:@19200.4]
  wire [15:0] _T_24281; // @[Mux.scala 19:72:@19201.4]
  wire [15:0] _T_24282; // @[Mux.scala 19:72:@19202.4]
  wire [15:0] _T_24283; // @[Mux.scala 19:72:@19203.4]
  wire [15:0] _T_24284; // @[Mux.scala 19:72:@19204.4]
  wire [15:0] _T_24285; // @[Mux.scala 19:72:@19205.4]
  wire [15:0] _T_24286; // @[Mux.scala 19:72:@19206.4]
  wire [15:0] _T_24287; // @[Mux.scala 19:72:@19207.4]
  wire [15:0] _T_24288; // @[Mux.scala 19:72:@19208.4]
  wire [15:0] _T_24289; // @[Mux.scala 19:72:@19209.4]
  wire [15:0] _T_24290; // @[Mux.scala 19:72:@19210.4]
  wire [15:0] _T_24291; // @[Mux.scala 19:72:@19211.4]
  wire [15:0] _T_24292; // @[Mux.scala 19:72:@19212.4]
  wire [15:0] _T_24293; // @[Mux.scala 19:72:@19213.4]
  wire [15:0] _T_24294; // @[Mux.scala 19:72:@19214.4]
  wire [7:0] _T_24872; // @[Mux.scala 19:72:@19564.4]
  wire [7:0] _T_24879; // @[Mux.scala 19:72:@19571.4]
  wire [15:0] _T_24880; // @[Mux.scala 19:72:@19572.4]
  wire [15:0] _T_24882; // @[Mux.scala 19:72:@19573.4]
  wire [7:0] _T_24889; // @[Mux.scala 19:72:@19580.4]
  wire [7:0] _T_24896; // @[Mux.scala 19:72:@19587.4]
  wire [15:0] _T_24897; // @[Mux.scala 19:72:@19588.4]
  wire [15:0] _T_24899; // @[Mux.scala 19:72:@19589.4]
  wire [7:0] _T_24906; // @[Mux.scala 19:72:@19596.4]
  wire [7:0] _T_24913; // @[Mux.scala 19:72:@19603.4]
  wire [15:0] _T_24914; // @[Mux.scala 19:72:@19604.4]
  wire [15:0] _T_24916; // @[Mux.scala 19:72:@19605.4]
  wire [7:0] _T_24923; // @[Mux.scala 19:72:@19612.4]
  wire [7:0] _T_24930; // @[Mux.scala 19:72:@19619.4]
  wire [15:0] _T_24931; // @[Mux.scala 19:72:@19620.4]
  wire [15:0] _T_24933; // @[Mux.scala 19:72:@19621.4]
  wire [7:0] _T_24940; // @[Mux.scala 19:72:@19628.4]
  wire [7:0] _T_24947; // @[Mux.scala 19:72:@19635.4]
  wire [15:0] _T_24948; // @[Mux.scala 19:72:@19636.4]
  wire [15:0] _T_24950; // @[Mux.scala 19:72:@19637.4]
  wire [7:0] _T_24957; // @[Mux.scala 19:72:@19644.4]
  wire [7:0] _T_24964; // @[Mux.scala 19:72:@19651.4]
  wire [15:0] _T_24965; // @[Mux.scala 19:72:@19652.4]
  wire [15:0] _T_24967; // @[Mux.scala 19:72:@19653.4]
  wire [7:0] _T_24974; // @[Mux.scala 19:72:@19660.4]
  wire [7:0] _T_24981; // @[Mux.scala 19:72:@19667.4]
  wire [15:0] _T_24982; // @[Mux.scala 19:72:@19668.4]
  wire [15:0] _T_24984; // @[Mux.scala 19:72:@19669.4]
  wire [7:0] _T_24991; // @[Mux.scala 19:72:@19676.4]
  wire [7:0] _T_24998; // @[Mux.scala 19:72:@19683.4]
  wire [15:0] _T_24999; // @[Mux.scala 19:72:@19684.4]
  wire [15:0] _T_25001; // @[Mux.scala 19:72:@19685.4]
  wire [15:0] _T_25016; // @[Mux.scala 19:72:@19700.4]
  wire [15:0] _T_25018; // @[Mux.scala 19:72:@19701.4]
  wire [15:0] _T_25033; // @[Mux.scala 19:72:@19716.4]
  wire [15:0] _T_25035; // @[Mux.scala 19:72:@19717.4]
  wire [15:0] _T_25050; // @[Mux.scala 19:72:@19732.4]
  wire [15:0] _T_25052; // @[Mux.scala 19:72:@19733.4]
  wire [15:0] _T_25067; // @[Mux.scala 19:72:@19748.4]
  wire [15:0] _T_25069; // @[Mux.scala 19:72:@19749.4]
  wire [15:0] _T_25084; // @[Mux.scala 19:72:@19764.4]
  wire [15:0] _T_25086; // @[Mux.scala 19:72:@19765.4]
  wire [15:0] _T_25101; // @[Mux.scala 19:72:@19780.4]
  wire [15:0] _T_25103; // @[Mux.scala 19:72:@19781.4]
  wire [15:0] _T_25118; // @[Mux.scala 19:72:@19796.4]
  wire [15:0] _T_25120; // @[Mux.scala 19:72:@19797.4]
  wire [15:0] _T_25135; // @[Mux.scala 19:72:@19812.4]
  wire [15:0] _T_25137; // @[Mux.scala 19:72:@19813.4]
  wire [15:0] _T_25138; // @[Mux.scala 19:72:@19814.4]
  wire [15:0] _T_25139; // @[Mux.scala 19:72:@19815.4]
  wire [15:0] _T_25140; // @[Mux.scala 19:72:@19816.4]
  wire [15:0] _T_25141; // @[Mux.scala 19:72:@19817.4]
  wire [15:0] _T_25142; // @[Mux.scala 19:72:@19818.4]
  wire [15:0] _T_25143; // @[Mux.scala 19:72:@19819.4]
  wire [15:0] _T_25144; // @[Mux.scala 19:72:@19820.4]
  wire [15:0] _T_25145; // @[Mux.scala 19:72:@19821.4]
  wire [15:0] _T_25146; // @[Mux.scala 19:72:@19822.4]
  wire [15:0] _T_25147; // @[Mux.scala 19:72:@19823.4]
  wire [15:0] _T_25148; // @[Mux.scala 19:72:@19824.4]
  wire [15:0] _T_25149; // @[Mux.scala 19:72:@19825.4]
  wire [15:0] _T_25150; // @[Mux.scala 19:72:@19826.4]
  wire [15:0] _T_25151; // @[Mux.scala 19:72:@19827.4]
  wire [15:0] _T_25152; // @[Mux.scala 19:72:@19828.4]
  wire [7:0] _T_25730; // @[Mux.scala 19:72:@20178.4]
  wire [7:0] _T_25737; // @[Mux.scala 19:72:@20185.4]
  wire [15:0] _T_25738; // @[Mux.scala 19:72:@20186.4]
  wire [15:0] _T_25740; // @[Mux.scala 19:72:@20187.4]
  wire [7:0] _T_25747; // @[Mux.scala 19:72:@20194.4]
  wire [7:0] _T_25754; // @[Mux.scala 19:72:@20201.4]
  wire [15:0] _T_25755; // @[Mux.scala 19:72:@20202.4]
  wire [15:0] _T_25757; // @[Mux.scala 19:72:@20203.4]
  wire [7:0] _T_25764; // @[Mux.scala 19:72:@20210.4]
  wire [7:0] _T_25771; // @[Mux.scala 19:72:@20217.4]
  wire [15:0] _T_25772; // @[Mux.scala 19:72:@20218.4]
  wire [15:0] _T_25774; // @[Mux.scala 19:72:@20219.4]
  wire [7:0] _T_25781; // @[Mux.scala 19:72:@20226.4]
  wire [7:0] _T_25788; // @[Mux.scala 19:72:@20233.4]
  wire [15:0] _T_25789; // @[Mux.scala 19:72:@20234.4]
  wire [15:0] _T_25791; // @[Mux.scala 19:72:@20235.4]
  wire [7:0] _T_25798; // @[Mux.scala 19:72:@20242.4]
  wire [7:0] _T_25805; // @[Mux.scala 19:72:@20249.4]
  wire [15:0] _T_25806; // @[Mux.scala 19:72:@20250.4]
  wire [15:0] _T_25808; // @[Mux.scala 19:72:@20251.4]
  wire [7:0] _T_25815; // @[Mux.scala 19:72:@20258.4]
  wire [7:0] _T_25822; // @[Mux.scala 19:72:@20265.4]
  wire [15:0] _T_25823; // @[Mux.scala 19:72:@20266.4]
  wire [15:0] _T_25825; // @[Mux.scala 19:72:@20267.4]
  wire [7:0] _T_25832; // @[Mux.scala 19:72:@20274.4]
  wire [7:0] _T_25839; // @[Mux.scala 19:72:@20281.4]
  wire [15:0] _T_25840; // @[Mux.scala 19:72:@20282.4]
  wire [15:0] _T_25842; // @[Mux.scala 19:72:@20283.4]
  wire [7:0] _T_25849; // @[Mux.scala 19:72:@20290.4]
  wire [7:0] _T_25856; // @[Mux.scala 19:72:@20297.4]
  wire [15:0] _T_25857; // @[Mux.scala 19:72:@20298.4]
  wire [15:0] _T_25859; // @[Mux.scala 19:72:@20299.4]
  wire [15:0] _T_25874; // @[Mux.scala 19:72:@20314.4]
  wire [15:0] _T_25876; // @[Mux.scala 19:72:@20315.4]
  wire [15:0] _T_25891; // @[Mux.scala 19:72:@20330.4]
  wire [15:0] _T_25893; // @[Mux.scala 19:72:@20331.4]
  wire [15:0] _T_25908; // @[Mux.scala 19:72:@20346.4]
  wire [15:0] _T_25910; // @[Mux.scala 19:72:@20347.4]
  wire [15:0] _T_25925; // @[Mux.scala 19:72:@20362.4]
  wire [15:0] _T_25927; // @[Mux.scala 19:72:@20363.4]
  wire [15:0] _T_25942; // @[Mux.scala 19:72:@20378.4]
  wire [15:0] _T_25944; // @[Mux.scala 19:72:@20379.4]
  wire [15:0] _T_25959; // @[Mux.scala 19:72:@20394.4]
  wire [15:0] _T_25961; // @[Mux.scala 19:72:@20395.4]
  wire [15:0] _T_25976; // @[Mux.scala 19:72:@20410.4]
  wire [15:0] _T_25978; // @[Mux.scala 19:72:@20411.4]
  wire [15:0] _T_25993; // @[Mux.scala 19:72:@20426.4]
  wire [15:0] _T_25995; // @[Mux.scala 19:72:@20427.4]
  wire [15:0] _T_25996; // @[Mux.scala 19:72:@20428.4]
  wire [15:0] _T_25997; // @[Mux.scala 19:72:@20429.4]
  wire [15:0] _T_25998; // @[Mux.scala 19:72:@20430.4]
  wire [15:0] _T_25999; // @[Mux.scala 19:72:@20431.4]
  wire [15:0] _T_26000; // @[Mux.scala 19:72:@20432.4]
  wire [15:0] _T_26001; // @[Mux.scala 19:72:@20433.4]
  wire [15:0] _T_26002; // @[Mux.scala 19:72:@20434.4]
  wire [15:0] _T_26003; // @[Mux.scala 19:72:@20435.4]
  wire [15:0] _T_26004; // @[Mux.scala 19:72:@20436.4]
  wire [15:0] _T_26005; // @[Mux.scala 19:72:@20437.4]
  wire [15:0] _T_26006; // @[Mux.scala 19:72:@20438.4]
  wire [15:0] _T_26007; // @[Mux.scala 19:72:@20439.4]
  wire [15:0] _T_26008; // @[Mux.scala 19:72:@20440.4]
  wire [15:0] _T_26009; // @[Mux.scala 19:72:@20441.4]
  wire [15:0] _T_26010; // @[Mux.scala 19:72:@20442.4]
  wire [7:0] _T_26588; // @[Mux.scala 19:72:@20792.4]
  wire [7:0] _T_26595; // @[Mux.scala 19:72:@20799.4]
  wire [15:0] _T_26596; // @[Mux.scala 19:72:@20800.4]
  wire [15:0] _T_26598; // @[Mux.scala 19:72:@20801.4]
  wire [7:0] _T_26605; // @[Mux.scala 19:72:@20808.4]
  wire [7:0] _T_26612; // @[Mux.scala 19:72:@20815.4]
  wire [15:0] _T_26613; // @[Mux.scala 19:72:@20816.4]
  wire [15:0] _T_26615; // @[Mux.scala 19:72:@20817.4]
  wire [7:0] _T_26622; // @[Mux.scala 19:72:@20824.4]
  wire [7:0] _T_26629; // @[Mux.scala 19:72:@20831.4]
  wire [15:0] _T_26630; // @[Mux.scala 19:72:@20832.4]
  wire [15:0] _T_26632; // @[Mux.scala 19:72:@20833.4]
  wire [7:0] _T_26639; // @[Mux.scala 19:72:@20840.4]
  wire [7:0] _T_26646; // @[Mux.scala 19:72:@20847.4]
  wire [15:0] _T_26647; // @[Mux.scala 19:72:@20848.4]
  wire [15:0] _T_26649; // @[Mux.scala 19:72:@20849.4]
  wire [7:0] _T_26656; // @[Mux.scala 19:72:@20856.4]
  wire [7:0] _T_26663; // @[Mux.scala 19:72:@20863.4]
  wire [15:0] _T_26664; // @[Mux.scala 19:72:@20864.4]
  wire [15:0] _T_26666; // @[Mux.scala 19:72:@20865.4]
  wire [7:0] _T_26673; // @[Mux.scala 19:72:@20872.4]
  wire [7:0] _T_26680; // @[Mux.scala 19:72:@20879.4]
  wire [15:0] _T_26681; // @[Mux.scala 19:72:@20880.4]
  wire [15:0] _T_26683; // @[Mux.scala 19:72:@20881.4]
  wire [7:0] _T_26690; // @[Mux.scala 19:72:@20888.4]
  wire [7:0] _T_26697; // @[Mux.scala 19:72:@20895.4]
  wire [15:0] _T_26698; // @[Mux.scala 19:72:@20896.4]
  wire [15:0] _T_26700; // @[Mux.scala 19:72:@20897.4]
  wire [7:0] _T_26707; // @[Mux.scala 19:72:@20904.4]
  wire [7:0] _T_26714; // @[Mux.scala 19:72:@20911.4]
  wire [15:0] _T_26715; // @[Mux.scala 19:72:@20912.4]
  wire [15:0] _T_26717; // @[Mux.scala 19:72:@20913.4]
  wire [15:0] _T_26732; // @[Mux.scala 19:72:@20928.4]
  wire [15:0] _T_26734; // @[Mux.scala 19:72:@20929.4]
  wire [15:0] _T_26749; // @[Mux.scala 19:72:@20944.4]
  wire [15:0] _T_26751; // @[Mux.scala 19:72:@20945.4]
  wire [15:0] _T_26766; // @[Mux.scala 19:72:@20960.4]
  wire [15:0] _T_26768; // @[Mux.scala 19:72:@20961.4]
  wire [15:0] _T_26783; // @[Mux.scala 19:72:@20976.4]
  wire [15:0] _T_26785; // @[Mux.scala 19:72:@20977.4]
  wire [15:0] _T_26800; // @[Mux.scala 19:72:@20992.4]
  wire [15:0] _T_26802; // @[Mux.scala 19:72:@20993.4]
  wire [15:0] _T_26817; // @[Mux.scala 19:72:@21008.4]
  wire [15:0] _T_26819; // @[Mux.scala 19:72:@21009.4]
  wire [15:0] _T_26834; // @[Mux.scala 19:72:@21024.4]
  wire [15:0] _T_26836; // @[Mux.scala 19:72:@21025.4]
  wire [15:0] _T_26851; // @[Mux.scala 19:72:@21040.4]
  wire [15:0] _T_26853; // @[Mux.scala 19:72:@21041.4]
  wire [15:0] _T_26854; // @[Mux.scala 19:72:@21042.4]
  wire [15:0] _T_26855; // @[Mux.scala 19:72:@21043.4]
  wire [15:0] _T_26856; // @[Mux.scala 19:72:@21044.4]
  wire [15:0] _T_26857; // @[Mux.scala 19:72:@21045.4]
  wire [15:0] _T_26858; // @[Mux.scala 19:72:@21046.4]
  wire [15:0] _T_26859; // @[Mux.scala 19:72:@21047.4]
  wire [15:0] _T_26860; // @[Mux.scala 19:72:@21048.4]
  wire [15:0] _T_26861; // @[Mux.scala 19:72:@21049.4]
  wire [15:0] _T_26862; // @[Mux.scala 19:72:@21050.4]
  wire [15:0] _T_26863; // @[Mux.scala 19:72:@21051.4]
  wire [15:0] _T_26864; // @[Mux.scala 19:72:@21052.4]
  wire [15:0] _T_26865; // @[Mux.scala 19:72:@21053.4]
  wire [15:0] _T_26866; // @[Mux.scala 19:72:@21054.4]
  wire [15:0] _T_26867; // @[Mux.scala 19:72:@21055.4]
  wire [15:0] _T_26868; // @[Mux.scala 19:72:@21056.4]
  wire [7:0] _T_27446; // @[Mux.scala 19:72:@21406.4]
  wire [7:0] _T_27453; // @[Mux.scala 19:72:@21413.4]
  wire [15:0] _T_27454; // @[Mux.scala 19:72:@21414.4]
  wire [15:0] _T_27456; // @[Mux.scala 19:72:@21415.4]
  wire [7:0] _T_27463; // @[Mux.scala 19:72:@21422.4]
  wire [7:0] _T_27470; // @[Mux.scala 19:72:@21429.4]
  wire [15:0] _T_27471; // @[Mux.scala 19:72:@21430.4]
  wire [15:0] _T_27473; // @[Mux.scala 19:72:@21431.4]
  wire [7:0] _T_27480; // @[Mux.scala 19:72:@21438.4]
  wire [7:0] _T_27487; // @[Mux.scala 19:72:@21445.4]
  wire [15:0] _T_27488; // @[Mux.scala 19:72:@21446.4]
  wire [15:0] _T_27490; // @[Mux.scala 19:72:@21447.4]
  wire [7:0] _T_27497; // @[Mux.scala 19:72:@21454.4]
  wire [7:0] _T_27504; // @[Mux.scala 19:72:@21461.4]
  wire [15:0] _T_27505; // @[Mux.scala 19:72:@21462.4]
  wire [15:0] _T_27507; // @[Mux.scala 19:72:@21463.4]
  wire [7:0] _T_27514; // @[Mux.scala 19:72:@21470.4]
  wire [7:0] _T_27521; // @[Mux.scala 19:72:@21477.4]
  wire [15:0] _T_27522; // @[Mux.scala 19:72:@21478.4]
  wire [15:0] _T_27524; // @[Mux.scala 19:72:@21479.4]
  wire [7:0] _T_27531; // @[Mux.scala 19:72:@21486.4]
  wire [7:0] _T_27538; // @[Mux.scala 19:72:@21493.4]
  wire [15:0] _T_27539; // @[Mux.scala 19:72:@21494.4]
  wire [15:0] _T_27541; // @[Mux.scala 19:72:@21495.4]
  wire [7:0] _T_27548; // @[Mux.scala 19:72:@21502.4]
  wire [7:0] _T_27555; // @[Mux.scala 19:72:@21509.4]
  wire [15:0] _T_27556; // @[Mux.scala 19:72:@21510.4]
  wire [15:0] _T_27558; // @[Mux.scala 19:72:@21511.4]
  wire [7:0] _T_27565; // @[Mux.scala 19:72:@21518.4]
  wire [7:0] _T_27572; // @[Mux.scala 19:72:@21525.4]
  wire [15:0] _T_27573; // @[Mux.scala 19:72:@21526.4]
  wire [15:0] _T_27575; // @[Mux.scala 19:72:@21527.4]
  wire [15:0] _T_27590; // @[Mux.scala 19:72:@21542.4]
  wire [15:0] _T_27592; // @[Mux.scala 19:72:@21543.4]
  wire [15:0] _T_27607; // @[Mux.scala 19:72:@21558.4]
  wire [15:0] _T_27609; // @[Mux.scala 19:72:@21559.4]
  wire [15:0] _T_27624; // @[Mux.scala 19:72:@21574.4]
  wire [15:0] _T_27626; // @[Mux.scala 19:72:@21575.4]
  wire [15:0] _T_27641; // @[Mux.scala 19:72:@21590.4]
  wire [15:0] _T_27643; // @[Mux.scala 19:72:@21591.4]
  wire [15:0] _T_27658; // @[Mux.scala 19:72:@21606.4]
  wire [15:0] _T_27660; // @[Mux.scala 19:72:@21607.4]
  wire [15:0] _T_27675; // @[Mux.scala 19:72:@21622.4]
  wire [15:0] _T_27677; // @[Mux.scala 19:72:@21623.4]
  wire [15:0] _T_27692; // @[Mux.scala 19:72:@21638.4]
  wire [15:0] _T_27694; // @[Mux.scala 19:72:@21639.4]
  wire [15:0] _T_27709; // @[Mux.scala 19:72:@21654.4]
  wire [15:0] _T_27711; // @[Mux.scala 19:72:@21655.4]
  wire [15:0] _T_27712; // @[Mux.scala 19:72:@21656.4]
  wire [15:0] _T_27713; // @[Mux.scala 19:72:@21657.4]
  wire [15:0] _T_27714; // @[Mux.scala 19:72:@21658.4]
  wire [15:0] _T_27715; // @[Mux.scala 19:72:@21659.4]
  wire [15:0] _T_27716; // @[Mux.scala 19:72:@21660.4]
  wire [15:0] _T_27717; // @[Mux.scala 19:72:@21661.4]
  wire [15:0] _T_27718; // @[Mux.scala 19:72:@21662.4]
  wire [15:0] _T_27719; // @[Mux.scala 19:72:@21663.4]
  wire [15:0] _T_27720; // @[Mux.scala 19:72:@21664.4]
  wire [15:0] _T_27721; // @[Mux.scala 19:72:@21665.4]
  wire [15:0] _T_27722; // @[Mux.scala 19:72:@21666.4]
  wire [15:0] _T_27723; // @[Mux.scala 19:72:@21667.4]
  wire [15:0] _T_27724; // @[Mux.scala 19:72:@21668.4]
  wire [15:0] _T_27725; // @[Mux.scala 19:72:@21669.4]
  wire [15:0] _T_27726; // @[Mux.scala 19:72:@21670.4]
  wire [7:0] _T_28304; // @[Mux.scala 19:72:@22020.4]
  wire [7:0] _T_28311; // @[Mux.scala 19:72:@22027.4]
  wire [15:0] _T_28312; // @[Mux.scala 19:72:@22028.4]
  wire [15:0] _T_28314; // @[Mux.scala 19:72:@22029.4]
  wire [7:0] _T_28321; // @[Mux.scala 19:72:@22036.4]
  wire [7:0] _T_28328; // @[Mux.scala 19:72:@22043.4]
  wire [15:0] _T_28329; // @[Mux.scala 19:72:@22044.4]
  wire [15:0] _T_28331; // @[Mux.scala 19:72:@22045.4]
  wire [7:0] _T_28338; // @[Mux.scala 19:72:@22052.4]
  wire [7:0] _T_28345; // @[Mux.scala 19:72:@22059.4]
  wire [15:0] _T_28346; // @[Mux.scala 19:72:@22060.4]
  wire [15:0] _T_28348; // @[Mux.scala 19:72:@22061.4]
  wire [7:0] _T_28355; // @[Mux.scala 19:72:@22068.4]
  wire [7:0] _T_28362; // @[Mux.scala 19:72:@22075.4]
  wire [15:0] _T_28363; // @[Mux.scala 19:72:@22076.4]
  wire [15:0] _T_28365; // @[Mux.scala 19:72:@22077.4]
  wire [7:0] _T_28372; // @[Mux.scala 19:72:@22084.4]
  wire [7:0] _T_28379; // @[Mux.scala 19:72:@22091.4]
  wire [15:0] _T_28380; // @[Mux.scala 19:72:@22092.4]
  wire [15:0] _T_28382; // @[Mux.scala 19:72:@22093.4]
  wire [7:0] _T_28389; // @[Mux.scala 19:72:@22100.4]
  wire [7:0] _T_28396; // @[Mux.scala 19:72:@22107.4]
  wire [15:0] _T_28397; // @[Mux.scala 19:72:@22108.4]
  wire [15:0] _T_28399; // @[Mux.scala 19:72:@22109.4]
  wire [7:0] _T_28406; // @[Mux.scala 19:72:@22116.4]
  wire [7:0] _T_28413; // @[Mux.scala 19:72:@22123.4]
  wire [15:0] _T_28414; // @[Mux.scala 19:72:@22124.4]
  wire [15:0] _T_28416; // @[Mux.scala 19:72:@22125.4]
  wire [7:0] _T_28423; // @[Mux.scala 19:72:@22132.4]
  wire [7:0] _T_28430; // @[Mux.scala 19:72:@22139.4]
  wire [15:0] _T_28431; // @[Mux.scala 19:72:@22140.4]
  wire [15:0] _T_28433; // @[Mux.scala 19:72:@22141.4]
  wire [15:0] _T_28448; // @[Mux.scala 19:72:@22156.4]
  wire [15:0] _T_28450; // @[Mux.scala 19:72:@22157.4]
  wire [15:0] _T_28465; // @[Mux.scala 19:72:@22172.4]
  wire [15:0] _T_28467; // @[Mux.scala 19:72:@22173.4]
  wire [15:0] _T_28482; // @[Mux.scala 19:72:@22188.4]
  wire [15:0] _T_28484; // @[Mux.scala 19:72:@22189.4]
  wire [15:0] _T_28499; // @[Mux.scala 19:72:@22204.4]
  wire [15:0] _T_28501; // @[Mux.scala 19:72:@22205.4]
  wire [15:0] _T_28516; // @[Mux.scala 19:72:@22220.4]
  wire [15:0] _T_28518; // @[Mux.scala 19:72:@22221.4]
  wire [15:0] _T_28533; // @[Mux.scala 19:72:@22236.4]
  wire [15:0] _T_28535; // @[Mux.scala 19:72:@22237.4]
  wire [15:0] _T_28550; // @[Mux.scala 19:72:@22252.4]
  wire [15:0] _T_28552; // @[Mux.scala 19:72:@22253.4]
  wire [15:0] _T_28567; // @[Mux.scala 19:72:@22268.4]
  wire [15:0] _T_28569; // @[Mux.scala 19:72:@22269.4]
  wire [15:0] _T_28570; // @[Mux.scala 19:72:@22270.4]
  wire [15:0] _T_28571; // @[Mux.scala 19:72:@22271.4]
  wire [15:0] _T_28572; // @[Mux.scala 19:72:@22272.4]
  wire [15:0] _T_28573; // @[Mux.scala 19:72:@22273.4]
  wire [15:0] _T_28574; // @[Mux.scala 19:72:@22274.4]
  wire [15:0] _T_28575; // @[Mux.scala 19:72:@22275.4]
  wire [15:0] _T_28576; // @[Mux.scala 19:72:@22276.4]
  wire [15:0] _T_28577; // @[Mux.scala 19:72:@22277.4]
  wire [15:0] _T_28578; // @[Mux.scala 19:72:@22278.4]
  wire [15:0] _T_28579; // @[Mux.scala 19:72:@22279.4]
  wire [15:0] _T_28580; // @[Mux.scala 19:72:@22280.4]
  wire [15:0] _T_28581; // @[Mux.scala 19:72:@22281.4]
  wire [15:0] _T_28582; // @[Mux.scala 19:72:@22282.4]
  wire [15:0] _T_28583; // @[Mux.scala 19:72:@22283.4]
  wire [15:0] _T_28584; // @[Mux.scala 19:72:@22284.4]
  wire [7:0] _T_29162; // @[Mux.scala 19:72:@22634.4]
  wire [7:0] _T_29169; // @[Mux.scala 19:72:@22641.4]
  wire [15:0] _T_29170; // @[Mux.scala 19:72:@22642.4]
  wire [15:0] _T_29172; // @[Mux.scala 19:72:@22643.4]
  wire [7:0] _T_29179; // @[Mux.scala 19:72:@22650.4]
  wire [7:0] _T_29186; // @[Mux.scala 19:72:@22657.4]
  wire [15:0] _T_29187; // @[Mux.scala 19:72:@22658.4]
  wire [15:0] _T_29189; // @[Mux.scala 19:72:@22659.4]
  wire [7:0] _T_29196; // @[Mux.scala 19:72:@22666.4]
  wire [7:0] _T_29203; // @[Mux.scala 19:72:@22673.4]
  wire [15:0] _T_29204; // @[Mux.scala 19:72:@22674.4]
  wire [15:0] _T_29206; // @[Mux.scala 19:72:@22675.4]
  wire [7:0] _T_29213; // @[Mux.scala 19:72:@22682.4]
  wire [7:0] _T_29220; // @[Mux.scala 19:72:@22689.4]
  wire [15:0] _T_29221; // @[Mux.scala 19:72:@22690.4]
  wire [15:0] _T_29223; // @[Mux.scala 19:72:@22691.4]
  wire [7:0] _T_29230; // @[Mux.scala 19:72:@22698.4]
  wire [7:0] _T_29237; // @[Mux.scala 19:72:@22705.4]
  wire [15:0] _T_29238; // @[Mux.scala 19:72:@22706.4]
  wire [15:0] _T_29240; // @[Mux.scala 19:72:@22707.4]
  wire [7:0] _T_29247; // @[Mux.scala 19:72:@22714.4]
  wire [7:0] _T_29254; // @[Mux.scala 19:72:@22721.4]
  wire [15:0] _T_29255; // @[Mux.scala 19:72:@22722.4]
  wire [15:0] _T_29257; // @[Mux.scala 19:72:@22723.4]
  wire [7:0] _T_29264; // @[Mux.scala 19:72:@22730.4]
  wire [7:0] _T_29271; // @[Mux.scala 19:72:@22737.4]
  wire [15:0] _T_29272; // @[Mux.scala 19:72:@22738.4]
  wire [15:0] _T_29274; // @[Mux.scala 19:72:@22739.4]
  wire [7:0] _T_29281; // @[Mux.scala 19:72:@22746.4]
  wire [7:0] _T_29288; // @[Mux.scala 19:72:@22753.4]
  wire [15:0] _T_29289; // @[Mux.scala 19:72:@22754.4]
  wire [15:0] _T_29291; // @[Mux.scala 19:72:@22755.4]
  wire [15:0] _T_29306; // @[Mux.scala 19:72:@22770.4]
  wire [15:0] _T_29308; // @[Mux.scala 19:72:@22771.4]
  wire [15:0] _T_29323; // @[Mux.scala 19:72:@22786.4]
  wire [15:0] _T_29325; // @[Mux.scala 19:72:@22787.4]
  wire [15:0] _T_29340; // @[Mux.scala 19:72:@22802.4]
  wire [15:0] _T_29342; // @[Mux.scala 19:72:@22803.4]
  wire [15:0] _T_29357; // @[Mux.scala 19:72:@22818.4]
  wire [15:0] _T_29359; // @[Mux.scala 19:72:@22819.4]
  wire [15:0] _T_29374; // @[Mux.scala 19:72:@22834.4]
  wire [15:0] _T_29376; // @[Mux.scala 19:72:@22835.4]
  wire [15:0] _T_29391; // @[Mux.scala 19:72:@22850.4]
  wire [15:0] _T_29393; // @[Mux.scala 19:72:@22851.4]
  wire [15:0] _T_29408; // @[Mux.scala 19:72:@22866.4]
  wire [15:0] _T_29410; // @[Mux.scala 19:72:@22867.4]
  wire [15:0] _T_29425; // @[Mux.scala 19:72:@22882.4]
  wire [15:0] _T_29427; // @[Mux.scala 19:72:@22883.4]
  wire [15:0] _T_29428; // @[Mux.scala 19:72:@22884.4]
  wire [15:0] _T_29429; // @[Mux.scala 19:72:@22885.4]
  wire [15:0] _T_29430; // @[Mux.scala 19:72:@22886.4]
  wire [15:0] _T_29431; // @[Mux.scala 19:72:@22887.4]
  wire [15:0] _T_29432; // @[Mux.scala 19:72:@22888.4]
  wire [15:0] _T_29433; // @[Mux.scala 19:72:@22889.4]
  wire [15:0] _T_29434; // @[Mux.scala 19:72:@22890.4]
  wire [15:0] _T_29435; // @[Mux.scala 19:72:@22891.4]
  wire [15:0] _T_29436; // @[Mux.scala 19:72:@22892.4]
  wire [15:0] _T_29437; // @[Mux.scala 19:72:@22893.4]
  wire [15:0] _T_29438; // @[Mux.scala 19:72:@22894.4]
  wire [15:0] _T_29439; // @[Mux.scala 19:72:@22895.4]
  wire [15:0] _T_29440; // @[Mux.scala 19:72:@22896.4]
  wire [15:0] _T_29441; // @[Mux.scala 19:72:@22897.4]
  wire [15:0] _T_29442; // @[Mux.scala 19:72:@22898.4]
  wire [7:0] _T_30020; // @[Mux.scala 19:72:@23248.4]
  wire [7:0] _T_30027; // @[Mux.scala 19:72:@23255.4]
  wire [15:0] _T_30028; // @[Mux.scala 19:72:@23256.4]
  wire [15:0] _T_30030; // @[Mux.scala 19:72:@23257.4]
  wire [7:0] _T_30037; // @[Mux.scala 19:72:@23264.4]
  wire [7:0] _T_30044; // @[Mux.scala 19:72:@23271.4]
  wire [15:0] _T_30045; // @[Mux.scala 19:72:@23272.4]
  wire [15:0] _T_30047; // @[Mux.scala 19:72:@23273.4]
  wire [7:0] _T_30054; // @[Mux.scala 19:72:@23280.4]
  wire [7:0] _T_30061; // @[Mux.scala 19:72:@23287.4]
  wire [15:0] _T_30062; // @[Mux.scala 19:72:@23288.4]
  wire [15:0] _T_30064; // @[Mux.scala 19:72:@23289.4]
  wire [7:0] _T_30071; // @[Mux.scala 19:72:@23296.4]
  wire [7:0] _T_30078; // @[Mux.scala 19:72:@23303.4]
  wire [15:0] _T_30079; // @[Mux.scala 19:72:@23304.4]
  wire [15:0] _T_30081; // @[Mux.scala 19:72:@23305.4]
  wire [7:0] _T_30088; // @[Mux.scala 19:72:@23312.4]
  wire [7:0] _T_30095; // @[Mux.scala 19:72:@23319.4]
  wire [15:0] _T_30096; // @[Mux.scala 19:72:@23320.4]
  wire [15:0] _T_30098; // @[Mux.scala 19:72:@23321.4]
  wire [7:0] _T_30105; // @[Mux.scala 19:72:@23328.4]
  wire [7:0] _T_30112; // @[Mux.scala 19:72:@23335.4]
  wire [15:0] _T_30113; // @[Mux.scala 19:72:@23336.4]
  wire [15:0] _T_30115; // @[Mux.scala 19:72:@23337.4]
  wire [7:0] _T_30122; // @[Mux.scala 19:72:@23344.4]
  wire [7:0] _T_30129; // @[Mux.scala 19:72:@23351.4]
  wire [15:0] _T_30130; // @[Mux.scala 19:72:@23352.4]
  wire [15:0] _T_30132; // @[Mux.scala 19:72:@23353.4]
  wire [7:0] _T_30139; // @[Mux.scala 19:72:@23360.4]
  wire [7:0] _T_30146; // @[Mux.scala 19:72:@23367.4]
  wire [15:0] _T_30147; // @[Mux.scala 19:72:@23368.4]
  wire [15:0] _T_30149; // @[Mux.scala 19:72:@23369.4]
  wire [15:0] _T_30164; // @[Mux.scala 19:72:@23384.4]
  wire [15:0] _T_30166; // @[Mux.scala 19:72:@23385.4]
  wire [15:0] _T_30181; // @[Mux.scala 19:72:@23400.4]
  wire [15:0] _T_30183; // @[Mux.scala 19:72:@23401.4]
  wire [15:0] _T_30198; // @[Mux.scala 19:72:@23416.4]
  wire [15:0] _T_30200; // @[Mux.scala 19:72:@23417.4]
  wire [15:0] _T_30215; // @[Mux.scala 19:72:@23432.4]
  wire [15:0] _T_30217; // @[Mux.scala 19:72:@23433.4]
  wire [15:0] _T_30232; // @[Mux.scala 19:72:@23448.4]
  wire [15:0] _T_30234; // @[Mux.scala 19:72:@23449.4]
  wire [15:0] _T_30249; // @[Mux.scala 19:72:@23464.4]
  wire [15:0] _T_30251; // @[Mux.scala 19:72:@23465.4]
  wire [15:0] _T_30266; // @[Mux.scala 19:72:@23480.4]
  wire [15:0] _T_30268; // @[Mux.scala 19:72:@23481.4]
  wire [15:0] _T_30283; // @[Mux.scala 19:72:@23496.4]
  wire [15:0] _T_30285; // @[Mux.scala 19:72:@23497.4]
  wire [15:0] _T_30286; // @[Mux.scala 19:72:@23498.4]
  wire [15:0] _T_30287; // @[Mux.scala 19:72:@23499.4]
  wire [15:0] _T_30288; // @[Mux.scala 19:72:@23500.4]
  wire [15:0] _T_30289; // @[Mux.scala 19:72:@23501.4]
  wire [15:0] _T_30290; // @[Mux.scala 19:72:@23502.4]
  wire [15:0] _T_30291; // @[Mux.scala 19:72:@23503.4]
  wire [15:0] _T_30292; // @[Mux.scala 19:72:@23504.4]
  wire [15:0] _T_30293; // @[Mux.scala 19:72:@23505.4]
  wire [15:0] _T_30294; // @[Mux.scala 19:72:@23506.4]
  wire [15:0] _T_30295; // @[Mux.scala 19:72:@23507.4]
  wire [15:0] _T_30296; // @[Mux.scala 19:72:@23508.4]
  wire [15:0] _T_30297; // @[Mux.scala 19:72:@23509.4]
  wire [15:0] _T_30298; // @[Mux.scala 19:72:@23510.4]
  wire [15:0] _T_30299; // @[Mux.scala 19:72:@23511.4]
  wire [15:0] _T_30300; // @[Mux.scala 19:72:@23512.4]
  wire [7:0] _T_30878; // @[Mux.scala 19:72:@23862.4]
  wire [7:0] _T_30885; // @[Mux.scala 19:72:@23869.4]
  wire [15:0] _T_30886; // @[Mux.scala 19:72:@23870.4]
  wire [15:0] _T_30888; // @[Mux.scala 19:72:@23871.4]
  wire [7:0] _T_30895; // @[Mux.scala 19:72:@23878.4]
  wire [7:0] _T_30902; // @[Mux.scala 19:72:@23885.4]
  wire [15:0] _T_30903; // @[Mux.scala 19:72:@23886.4]
  wire [15:0] _T_30905; // @[Mux.scala 19:72:@23887.4]
  wire [7:0] _T_30912; // @[Mux.scala 19:72:@23894.4]
  wire [7:0] _T_30919; // @[Mux.scala 19:72:@23901.4]
  wire [15:0] _T_30920; // @[Mux.scala 19:72:@23902.4]
  wire [15:0] _T_30922; // @[Mux.scala 19:72:@23903.4]
  wire [7:0] _T_30929; // @[Mux.scala 19:72:@23910.4]
  wire [7:0] _T_30936; // @[Mux.scala 19:72:@23917.4]
  wire [15:0] _T_30937; // @[Mux.scala 19:72:@23918.4]
  wire [15:0] _T_30939; // @[Mux.scala 19:72:@23919.4]
  wire [7:0] _T_30946; // @[Mux.scala 19:72:@23926.4]
  wire [7:0] _T_30953; // @[Mux.scala 19:72:@23933.4]
  wire [15:0] _T_30954; // @[Mux.scala 19:72:@23934.4]
  wire [15:0] _T_30956; // @[Mux.scala 19:72:@23935.4]
  wire [7:0] _T_30963; // @[Mux.scala 19:72:@23942.4]
  wire [7:0] _T_30970; // @[Mux.scala 19:72:@23949.4]
  wire [15:0] _T_30971; // @[Mux.scala 19:72:@23950.4]
  wire [15:0] _T_30973; // @[Mux.scala 19:72:@23951.4]
  wire [7:0] _T_30980; // @[Mux.scala 19:72:@23958.4]
  wire [7:0] _T_30987; // @[Mux.scala 19:72:@23965.4]
  wire [15:0] _T_30988; // @[Mux.scala 19:72:@23966.4]
  wire [15:0] _T_30990; // @[Mux.scala 19:72:@23967.4]
  wire [7:0] _T_30997; // @[Mux.scala 19:72:@23974.4]
  wire [7:0] _T_31004; // @[Mux.scala 19:72:@23981.4]
  wire [15:0] _T_31005; // @[Mux.scala 19:72:@23982.4]
  wire [15:0] _T_31007; // @[Mux.scala 19:72:@23983.4]
  wire [15:0] _T_31022; // @[Mux.scala 19:72:@23998.4]
  wire [15:0] _T_31024; // @[Mux.scala 19:72:@23999.4]
  wire [15:0] _T_31039; // @[Mux.scala 19:72:@24014.4]
  wire [15:0] _T_31041; // @[Mux.scala 19:72:@24015.4]
  wire [15:0] _T_31056; // @[Mux.scala 19:72:@24030.4]
  wire [15:0] _T_31058; // @[Mux.scala 19:72:@24031.4]
  wire [15:0] _T_31073; // @[Mux.scala 19:72:@24046.4]
  wire [15:0] _T_31075; // @[Mux.scala 19:72:@24047.4]
  wire [15:0] _T_31090; // @[Mux.scala 19:72:@24062.4]
  wire [15:0] _T_31092; // @[Mux.scala 19:72:@24063.4]
  wire [15:0] _T_31107; // @[Mux.scala 19:72:@24078.4]
  wire [15:0] _T_31109; // @[Mux.scala 19:72:@24079.4]
  wire [15:0] _T_31124; // @[Mux.scala 19:72:@24094.4]
  wire [15:0] _T_31126; // @[Mux.scala 19:72:@24095.4]
  wire [15:0] _T_31141; // @[Mux.scala 19:72:@24110.4]
  wire [15:0] _T_31143; // @[Mux.scala 19:72:@24111.4]
  wire [15:0] _T_31144; // @[Mux.scala 19:72:@24112.4]
  wire [15:0] _T_31145; // @[Mux.scala 19:72:@24113.4]
  wire [15:0] _T_31146; // @[Mux.scala 19:72:@24114.4]
  wire [15:0] _T_31147; // @[Mux.scala 19:72:@24115.4]
  wire [15:0] _T_31148; // @[Mux.scala 19:72:@24116.4]
  wire [15:0] _T_31149; // @[Mux.scala 19:72:@24117.4]
  wire [15:0] _T_31150; // @[Mux.scala 19:72:@24118.4]
  wire [15:0] _T_31151; // @[Mux.scala 19:72:@24119.4]
  wire [15:0] _T_31152; // @[Mux.scala 19:72:@24120.4]
  wire [15:0] _T_31153; // @[Mux.scala 19:72:@24121.4]
  wire [15:0] _T_31154; // @[Mux.scala 19:72:@24122.4]
  wire [15:0] _T_31155; // @[Mux.scala 19:72:@24123.4]
  wire [15:0] _T_31156; // @[Mux.scala 19:72:@24124.4]
  wire [15:0] _T_31157; // @[Mux.scala 19:72:@24125.4]
  wire [15:0] _T_31158; // @[Mux.scala 19:72:@24126.4]
  reg  conflictPReg_0_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_163;
  reg  conflictPReg_0_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_164;
  reg  conflictPReg_0_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_165;
  reg  conflictPReg_0_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_166;
  reg  conflictPReg_0_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_167;
  reg  conflictPReg_0_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_168;
  reg  conflictPReg_0_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_169;
  reg  conflictPReg_0_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_170;
  reg  conflictPReg_0_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_171;
  reg  conflictPReg_0_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_172;
  reg  conflictPReg_0_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_173;
  reg  conflictPReg_0_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_174;
  reg  conflictPReg_0_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_175;
  reg  conflictPReg_0_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_176;
  reg  conflictPReg_0_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_177;
  reg  conflictPReg_0_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_178;
  reg  conflictPReg_1_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_179;
  reg  conflictPReg_1_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_180;
  reg  conflictPReg_1_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_181;
  reg  conflictPReg_1_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_182;
  reg  conflictPReg_1_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_183;
  reg  conflictPReg_1_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_184;
  reg  conflictPReg_1_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_185;
  reg  conflictPReg_1_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_186;
  reg  conflictPReg_1_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_187;
  reg  conflictPReg_1_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_188;
  reg  conflictPReg_1_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_189;
  reg  conflictPReg_1_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_190;
  reg  conflictPReg_1_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_191;
  reg  conflictPReg_1_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_192;
  reg  conflictPReg_1_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_193;
  reg  conflictPReg_1_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_194;
  reg  conflictPReg_2_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_195;
  reg  conflictPReg_2_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_196;
  reg  conflictPReg_2_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_197;
  reg  conflictPReg_2_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_198;
  reg  conflictPReg_2_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_199;
  reg  conflictPReg_2_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_200;
  reg  conflictPReg_2_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_201;
  reg  conflictPReg_2_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_202;
  reg  conflictPReg_2_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_203;
  reg  conflictPReg_2_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_204;
  reg  conflictPReg_2_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_205;
  reg  conflictPReg_2_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_206;
  reg  conflictPReg_2_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_207;
  reg  conflictPReg_2_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_208;
  reg  conflictPReg_2_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_209;
  reg  conflictPReg_2_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_210;
  reg  conflictPReg_3_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_211;
  reg  conflictPReg_3_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_212;
  reg  conflictPReg_3_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_213;
  reg  conflictPReg_3_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_214;
  reg  conflictPReg_3_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_215;
  reg  conflictPReg_3_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_216;
  reg  conflictPReg_3_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_217;
  reg  conflictPReg_3_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_218;
  reg  conflictPReg_3_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_219;
  reg  conflictPReg_3_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_220;
  reg  conflictPReg_3_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_221;
  reg  conflictPReg_3_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_222;
  reg  conflictPReg_3_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_223;
  reg  conflictPReg_3_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_224;
  reg  conflictPReg_3_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_225;
  reg  conflictPReg_3_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_226;
  reg  conflictPReg_4_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_227;
  reg  conflictPReg_4_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_228;
  reg  conflictPReg_4_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_229;
  reg  conflictPReg_4_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_230;
  reg  conflictPReg_4_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_231;
  reg  conflictPReg_4_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_232;
  reg  conflictPReg_4_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_233;
  reg  conflictPReg_4_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_234;
  reg  conflictPReg_4_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_235;
  reg  conflictPReg_4_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_236;
  reg  conflictPReg_4_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_237;
  reg  conflictPReg_4_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_238;
  reg  conflictPReg_4_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_239;
  reg  conflictPReg_4_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_240;
  reg  conflictPReg_4_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_241;
  reg  conflictPReg_4_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_242;
  reg  conflictPReg_5_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_243;
  reg  conflictPReg_5_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_244;
  reg  conflictPReg_5_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_245;
  reg  conflictPReg_5_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_246;
  reg  conflictPReg_5_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_247;
  reg  conflictPReg_5_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_248;
  reg  conflictPReg_5_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_249;
  reg  conflictPReg_5_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_250;
  reg  conflictPReg_5_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_251;
  reg  conflictPReg_5_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_252;
  reg  conflictPReg_5_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_253;
  reg  conflictPReg_5_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_254;
  reg  conflictPReg_5_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_255;
  reg  conflictPReg_5_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_256;
  reg  conflictPReg_5_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_257;
  reg  conflictPReg_5_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_258;
  reg  conflictPReg_6_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_259;
  reg  conflictPReg_6_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_260;
  reg  conflictPReg_6_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_261;
  reg  conflictPReg_6_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_262;
  reg  conflictPReg_6_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_263;
  reg  conflictPReg_6_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_264;
  reg  conflictPReg_6_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_265;
  reg  conflictPReg_6_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_266;
  reg  conflictPReg_6_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_267;
  reg  conflictPReg_6_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_268;
  reg  conflictPReg_6_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_269;
  reg  conflictPReg_6_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_270;
  reg  conflictPReg_6_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_271;
  reg  conflictPReg_6_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_272;
  reg  conflictPReg_6_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_273;
  reg  conflictPReg_6_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_274;
  reg  conflictPReg_7_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_275;
  reg  conflictPReg_7_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_276;
  reg  conflictPReg_7_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_277;
  reg  conflictPReg_7_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_278;
  reg  conflictPReg_7_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_279;
  reg  conflictPReg_7_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_280;
  reg  conflictPReg_7_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_281;
  reg  conflictPReg_7_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_282;
  reg  conflictPReg_7_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_283;
  reg  conflictPReg_7_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_284;
  reg  conflictPReg_7_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_285;
  reg  conflictPReg_7_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_286;
  reg  conflictPReg_7_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_287;
  reg  conflictPReg_7_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_288;
  reg  conflictPReg_7_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_289;
  reg  conflictPReg_7_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_290;
  reg  conflictPReg_8_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_291;
  reg  conflictPReg_8_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_292;
  reg  conflictPReg_8_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_293;
  reg  conflictPReg_8_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_294;
  reg  conflictPReg_8_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_295;
  reg  conflictPReg_8_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_296;
  reg  conflictPReg_8_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_297;
  reg  conflictPReg_8_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_298;
  reg  conflictPReg_8_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_299;
  reg  conflictPReg_8_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_300;
  reg  conflictPReg_8_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_301;
  reg  conflictPReg_8_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_302;
  reg  conflictPReg_8_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_303;
  reg  conflictPReg_8_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_304;
  reg  conflictPReg_8_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_305;
  reg  conflictPReg_8_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_306;
  reg  conflictPReg_9_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_307;
  reg  conflictPReg_9_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_308;
  reg  conflictPReg_9_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_309;
  reg  conflictPReg_9_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_310;
  reg  conflictPReg_9_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_311;
  reg  conflictPReg_9_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_312;
  reg  conflictPReg_9_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_313;
  reg  conflictPReg_9_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_314;
  reg  conflictPReg_9_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_315;
  reg  conflictPReg_9_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_316;
  reg  conflictPReg_9_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_317;
  reg  conflictPReg_9_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_318;
  reg  conflictPReg_9_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_319;
  reg  conflictPReg_9_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_320;
  reg  conflictPReg_9_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_321;
  reg  conflictPReg_9_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_322;
  reg  conflictPReg_10_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_323;
  reg  conflictPReg_10_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_324;
  reg  conflictPReg_10_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_325;
  reg  conflictPReg_10_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_326;
  reg  conflictPReg_10_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_327;
  reg  conflictPReg_10_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_328;
  reg  conflictPReg_10_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_329;
  reg  conflictPReg_10_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_330;
  reg  conflictPReg_10_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_331;
  reg  conflictPReg_10_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_332;
  reg  conflictPReg_10_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_333;
  reg  conflictPReg_10_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_334;
  reg  conflictPReg_10_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_335;
  reg  conflictPReg_10_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_336;
  reg  conflictPReg_10_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_337;
  reg  conflictPReg_10_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_338;
  reg  conflictPReg_11_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_339;
  reg  conflictPReg_11_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_340;
  reg  conflictPReg_11_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_341;
  reg  conflictPReg_11_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_342;
  reg  conflictPReg_11_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_343;
  reg  conflictPReg_11_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_344;
  reg  conflictPReg_11_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_345;
  reg  conflictPReg_11_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_346;
  reg  conflictPReg_11_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_347;
  reg  conflictPReg_11_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_348;
  reg  conflictPReg_11_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_349;
  reg  conflictPReg_11_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_350;
  reg  conflictPReg_11_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_351;
  reg  conflictPReg_11_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_352;
  reg  conflictPReg_11_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_353;
  reg  conflictPReg_11_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_354;
  reg  conflictPReg_12_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_355;
  reg  conflictPReg_12_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_356;
  reg  conflictPReg_12_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_357;
  reg  conflictPReg_12_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_358;
  reg  conflictPReg_12_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_359;
  reg  conflictPReg_12_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_360;
  reg  conflictPReg_12_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_361;
  reg  conflictPReg_12_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_362;
  reg  conflictPReg_12_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_363;
  reg  conflictPReg_12_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_364;
  reg  conflictPReg_12_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_365;
  reg  conflictPReg_12_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_366;
  reg  conflictPReg_12_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_367;
  reg  conflictPReg_12_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_368;
  reg  conflictPReg_12_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_369;
  reg  conflictPReg_12_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_370;
  reg  conflictPReg_13_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_371;
  reg  conflictPReg_13_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_372;
  reg  conflictPReg_13_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_373;
  reg  conflictPReg_13_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_374;
  reg  conflictPReg_13_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_375;
  reg  conflictPReg_13_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_376;
  reg  conflictPReg_13_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_377;
  reg  conflictPReg_13_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_378;
  reg  conflictPReg_13_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_379;
  reg  conflictPReg_13_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_380;
  reg  conflictPReg_13_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_381;
  reg  conflictPReg_13_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_382;
  reg  conflictPReg_13_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_383;
  reg  conflictPReg_13_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_384;
  reg  conflictPReg_13_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_385;
  reg  conflictPReg_13_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_386;
  reg  conflictPReg_14_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_387;
  reg  conflictPReg_14_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_388;
  reg  conflictPReg_14_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_389;
  reg  conflictPReg_14_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_390;
  reg  conflictPReg_14_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_391;
  reg  conflictPReg_14_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_392;
  reg  conflictPReg_14_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_393;
  reg  conflictPReg_14_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_394;
  reg  conflictPReg_14_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_395;
  reg  conflictPReg_14_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_396;
  reg  conflictPReg_14_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_397;
  reg  conflictPReg_14_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_398;
  reg  conflictPReg_14_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_399;
  reg  conflictPReg_14_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_400;
  reg  conflictPReg_14_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_401;
  reg  conflictPReg_14_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_402;
  reg  conflictPReg_15_0; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_403;
  reg  conflictPReg_15_1; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_404;
  reg  conflictPReg_15_2; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_405;
  reg  conflictPReg_15_3; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_406;
  reg  conflictPReg_15_4; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_407;
  reg  conflictPReg_15_5; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_408;
  reg  conflictPReg_15_6; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_409;
  reg  conflictPReg_15_7; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_410;
  reg  conflictPReg_15_8; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_411;
  reg  conflictPReg_15_9; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_412;
  reg  conflictPReg_15_10; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_413;
  reg  conflictPReg_15_11; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_414;
  reg  conflictPReg_15_12; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_415;
  reg  conflictPReg_15_13; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_416;
  reg  conflictPReg_15_14; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_417;
  reg  conflictPReg_15_15; // @[AxiLoadQueue.scala 166:29:@24419.4]
  reg [31:0] _RAND_418;
  wire [7:0] _T_52332; // @[Mux.scala 19:72:@24990.4]
  wire [7:0] _T_52339; // @[Mux.scala 19:72:@24997.4]
  wire [15:0] _T_52340; // @[Mux.scala 19:72:@24998.4]
  wire [15:0] _T_52342; // @[Mux.scala 19:72:@24999.4]
  wire [7:0] _T_52349; // @[Mux.scala 19:72:@25006.4]
  wire [7:0] _T_52356; // @[Mux.scala 19:72:@25013.4]
  wire [15:0] _T_52357; // @[Mux.scala 19:72:@25014.4]
  wire [15:0] _T_52359; // @[Mux.scala 19:72:@25015.4]
  wire [7:0] _T_52366; // @[Mux.scala 19:72:@25022.4]
  wire [7:0] _T_52373; // @[Mux.scala 19:72:@25029.4]
  wire [15:0] _T_52374; // @[Mux.scala 19:72:@25030.4]
  wire [15:0] _T_52376; // @[Mux.scala 19:72:@25031.4]
  wire [7:0] _T_52383; // @[Mux.scala 19:72:@25038.4]
  wire [7:0] _T_52390; // @[Mux.scala 19:72:@25045.4]
  wire [15:0] _T_52391; // @[Mux.scala 19:72:@25046.4]
  wire [15:0] _T_52393; // @[Mux.scala 19:72:@25047.4]
  wire [7:0] _T_52400; // @[Mux.scala 19:72:@25054.4]
  wire [7:0] _T_52407; // @[Mux.scala 19:72:@25061.4]
  wire [15:0] _T_52408; // @[Mux.scala 19:72:@25062.4]
  wire [15:0] _T_52410; // @[Mux.scala 19:72:@25063.4]
  wire [7:0] _T_52417; // @[Mux.scala 19:72:@25070.4]
  wire [7:0] _T_52424; // @[Mux.scala 19:72:@25077.4]
  wire [15:0] _T_52425; // @[Mux.scala 19:72:@25078.4]
  wire [15:0] _T_52427; // @[Mux.scala 19:72:@25079.4]
  wire [7:0] _T_52434; // @[Mux.scala 19:72:@25086.4]
  wire [7:0] _T_52441; // @[Mux.scala 19:72:@25093.4]
  wire [15:0] _T_52442; // @[Mux.scala 19:72:@25094.4]
  wire [15:0] _T_52444; // @[Mux.scala 19:72:@25095.4]
  wire [7:0] _T_52451; // @[Mux.scala 19:72:@25102.4]
  wire [7:0] _T_52458; // @[Mux.scala 19:72:@25109.4]
  wire [15:0] _T_52459; // @[Mux.scala 19:72:@25110.4]
  wire [15:0] _T_52461; // @[Mux.scala 19:72:@25111.4]
  wire [15:0] _T_52476; // @[Mux.scala 19:72:@25126.4]
  wire [15:0] _T_52478; // @[Mux.scala 19:72:@25127.4]
  wire [15:0] _T_52493; // @[Mux.scala 19:72:@25142.4]
  wire [15:0] _T_52495; // @[Mux.scala 19:72:@25143.4]
  wire [15:0] _T_52510; // @[Mux.scala 19:72:@25158.4]
  wire [15:0] _T_52512; // @[Mux.scala 19:72:@25159.4]
  wire [15:0] _T_52527; // @[Mux.scala 19:72:@25174.4]
  wire [15:0] _T_52529; // @[Mux.scala 19:72:@25175.4]
  wire [15:0] _T_52544; // @[Mux.scala 19:72:@25190.4]
  wire [15:0] _T_52546; // @[Mux.scala 19:72:@25191.4]
  wire [15:0] _T_52561; // @[Mux.scala 19:72:@25206.4]
  wire [15:0] _T_52563; // @[Mux.scala 19:72:@25207.4]
  wire [15:0] _T_52578; // @[Mux.scala 19:72:@25222.4]
  wire [15:0] _T_52580; // @[Mux.scala 19:72:@25223.4]
  wire [15:0] _T_52595; // @[Mux.scala 19:72:@25238.4]
  wire [15:0] _T_52597; // @[Mux.scala 19:72:@25239.4]
  wire [15:0] _T_52598; // @[Mux.scala 19:72:@25240.4]
  wire [15:0] _T_52599; // @[Mux.scala 19:72:@25241.4]
  wire [15:0] _T_52600; // @[Mux.scala 19:72:@25242.4]
  wire [15:0] _T_52601; // @[Mux.scala 19:72:@25243.4]
  wire [15:0] _T_52602; // @[Mux.scala 19:72:@25244.4]
  wire [15:0] _T_52603; // @[Mux.scala 19:72:@25245.4]
  wire [15:0] _T_52604; // @[Mux.scala 19:72:@25246.4]
  wire [15:0] _T_52605; // @[Mux.scala 19:72:@25247.4]
  wire [15:0] _T_52606; // @[Mux.scala 19:72:@25248.4]
  wire [15:0] _T_52607; // @[Mux.scala 19:72:@25249.4]
  wire [15:0] _T_52608; // @[Mux.scala 19:72:@25250.4]
  wire [15:0] _T_52609; // @[Mux.scala 19:72:@25251.4]
  wire [15:0] _T_52610; // @[Mux.scala 19:72:@25252.4]
  wire [15:0] _T_52611; // @[Mux.scala 19:72:@25253.4]
  wire [15:0] _T_52612; // @[Mux.scala 19:72:@25254.4]
  wire [7:0] _T_53190; // @[Mux.scala 19:72:@25604.4]
  wire [7:0] _T_53197; // @[Mux.scala 19:72:@25611.4]
  wire [15:0] _T_53198; // @[Mux.scala 19:72:@25612.4]
  wire [15:0] _T_53200; // @[Mux.scala 19:72:@25613.4]
  wire [7:0] _T_53207; // @[Mux.scala 19:72:@25620.4]
  wire [7:0] _T_53214; // @[Mux.scala 19:72:@25627.4]
  wire [15:0] _T_53215; // @[Mux.scala 19:72:@25628.4]
  wire [15:0] _T_53217; // @[Mux.scala 19:72:@25629.4]
  wire [7:0] _T_53224; // @[Mux.scala 19:72:@25636.4]
  wire [7:0] _T_53231; // @[Mux.scala 19:72:@25643.4]
  wire [15:0] _T_53232; // @[Mux.scala 19:72:@25644.4]
  wire [15:0] _T_53234; // @[Mux.scala 19:72:@25645.4]
  wire [7:0] _T_53241; // @[Mux.scala 19:72:@25652.4]
  wire [7:0] _T_53248; // @[Mux.scala 19:72:@25659.4]
  wire [15:0] _T_53249; // @[Mux.scala 19:72:@25660.4]
  wire [15:0] _T_53251; // @[Mux.scala 19:72:@25661.4]
  wire [7:0] _T_53258; // @[Mux.scala 19:72:@25668.4]
  wire [7:0] _T_53265; // @[Mux.scala 19:72:@25675.4]
  wire [15:0] _T_53266; // @[Mux.scala 19:72:@25676.4]
  wire [15:0] _T_53268; // @[Mux.scala 19:72:@25677.4]
  wire [7:0] _T_53275; // @[Mux.scala 19:72:@25684.4]
  wire [7:0] _T_53282; // @[Mux.scala 19:72:@25691.4]
  wire [15:0] _T_53283; // @[Mux.scala 19:72:@25692.4]
  wire [15:0] _T_53285; // @[Mux.scala 19:72:@25693.4]
  wire [7:0] _T_53292; // @[Mux.scala 19:72:@25700.4]
  wire [7:0] _T_53299; // @[Mux.scala 19:72:@25707.4]
  wire [15:0] _T_53300; // @[Mux.scala 19:72:@25708.4]
  wire [15:0] _T_53302; // @[Mux.scala 19:72:@25709.4]
  wire [7:0] _T_53309; // @[Mux.scala 19:72:@25716.4]
  wire [7:0] _T_53316; // @[Mux.scala 19:72:@25723.4]
  wire [15:0] _T_53317; // @[Mux.scala 19:72:@25724.4]
  wire [15:0] _T_53319; // @[Mux.scala 19:72:@25725.4]
  wire [15:0] _T_53334; // @[Mux.scala 19:72:@25740.4]
  wire [15:0] _T_53336; // @[Mux.scala 19:72:@25741.4]
  wire [15:0] _T_53351; // @[Mux.scala 19:72:@25756.4]
  wire [15:0] _T_53353; // @[Mux.scala 19:72:@25757.4]
  wire [15:0] _T_53368; // @[Mux.scala 19:72:@25772.4]
  wire [15:0] _T_53370; // @[Mux.scala 19:72:@25773.4]
  wire [15:0] _T_53385; // @[Mux.scala 19:72:@25788.4]
  wire [15:0] _T_53387; // @[Mux.scala 19:72:@25789.4]
  wire [15:0] _T_53402; // @[Mux.scala 19:72:@25804.4]
  wire [15:0] _T_53404; // @[Mux.scala 19:72:@25805.4]
  wire [15:0] _T_53419; // @[Mux.scala 19:72:@25820.4]
  wire [15:0] _T_53421; // @[Mux.scala 19:72:@25821.4]
  wire [15:0] _T_53436; // @[Mux.scala 19:72:@25836.4]
  wire [15:0] _T_53438; // @[Mux.scala 19:72:@25837.4]
  wire [15:0] _T_53453; // @[Mux.scala 19:72:@25852.4]
  wire [15:0] _T_53455; // @[Mux.scala 19:72:@25853.4]
  wire [15:0] _T_53456; // @[Mux.scala 19:72:@25854.4]
  wire [15:0] _T_53457; // @[Mux.scala 19:72:@25855.4]
  wire [15:0] _T_53458; // @[Mux.scala 19:72:@25856.4]
  wire [15:0] _T_53459; // @[Mux.scala 19:72:@25857.4]
  wire [15:0] _T_53460; // @[Mux.scala 19:72:@25858.4]
  wire [15:0] _T_53461; // @[Mux.scala 19:72:@25859.4]
  wire [15:0] _T_53462; // @[Mux.scala 19:72:@25860.4]
  wire [15:0] _T_53463; // @[Mux.scala 19:72:@25861.4]
  wire [15:0] _T_53464; // @[Mux.scala 19:72:@25862.4]
  wire [15:0] _T_53465; // @[Mux.scala 19:72:@25863.4]
  wire [15:0] _T_53466; // @[Mux.scala 19:72:@25864.4]
  wire [15:0] _T_53467; // @[Mux.scala 19:72:@25865.4]
  wire [15:0] _T_53468; // @[Mux.scala 19:72:@25866.4]
  wire [15:0] _T_53469; // @[Mux.scala 19:72:@25867.4]
  wire [15:0] _T_53470; // @[Mux.scala 19:72:@25868.4]
  wire [7:0] _T_54048; // @[Mux.scala 19:72:@26218.4]
  wire [7:0] _T_54055; // @[Mux.scala 19:72:@26225.4]
  wire [15:0] _T_54056; // @[Mux.scala 19:72:@26226.4]
  wire [15:0] _T_54058; // @[Mux.scala 19:72:@26227.4]
  wire [7:0] _T_54065; // @[Mux.scala 19:72:@26234.4]
  wire [7:0] _T_54072; // @[Mux.scala 19:72:@26241.4]
  wire [15:0] _T_54073; // @[Mux.scala 19:72:@26242.4]
  wire [15:0] _T_54075; // @[Mux.scala 19:72:@26243.4]
  wire [7:0] _T_54082; // @[Mux.scala 19:72:@26250.4]
  wire [7:0] _T_54089; // @[Mux.scala 19:72:@26257.4]
  wire [15:0] _T_54090; // @[Mux.scala 19:72:@26258.4]
  wire [15:0] _T_54092; // @[Mux.scala 19:72:@26259.4]
  wire [7:0] _T_54099; // @[Mux.scala 19:72:@26266.4]
  wire [7:0] _T_54106; // @[Mux.scala 19:72:@26273.4]
  wire [15:0] _T_54107; // @[Mux.scala 19:72:@26274.4]
  wire [15:0] _T_54109; // @[Mux.scala 19:72:@26275.4]
  wire [7:0] _T_54116; // @[Mux.scala 19:72:@26282.4]
  wire [7:0] _T_54123; // @[Mux.scala 19:72:@26289.4]
  wire [15:0] _T_54124; // @[Mux.scala 19:72:@26290.4]
  wire [15:0] _T_54126; // @[Mux.scala 19:72:@26291.4]
  wire [7:0] _T_54133; // @[Mux.scala 19:72:@26298.4]
  wire [7:0] _T_54140; // @[Mux.scala 19:72:@26305.4]
  wire [15:0] _T_54141; // @[Mux.scala 19:72:@26306.4]
  wire [15:0] _T_54143; // @[Mux.scala 19:72:@26307.4]
  wire [7:0] _T_54150; // @[Mux.scala 19:72:@26314.4]
  wire [7:0] _T_54157; // @[Mux.scala 19:72:@26321.4]
  wire [15:0] _T_54158; // @[Mux.scala 19:72:@26322.4]
  wire [15:0] _T_54160; // @[Mux.scala 19:72:@26323.4]
  wire [7:0] _T_54167; // @[Mux.scala 19:72:@26330.4]
  wire [7:0] _T_54174; // @[Mux.scala 19:72:@26337.4]
  wire [15:0] _T_54175; // @[Mux.scala 19:72:@26338.4]
  wire [15:0] _T_54177; // @[Mux.scala 19:72:@26339.4]
  wire [15:0] _T_54192; // @[Mux.scala 19:72:@26354.4]
  wire [15:0] _T_54194; // @[Mux.scala 19:72:@26355.4]
  wire [15:0] _T_54209; // @[Mux.scala 19:72:@26370.4]
  wire [15:0] _T_54211; // @[Mux.scala 19:72:@26371.4]
  wire [15:0] _T_54226; // @[Mux.scala 19:72:@26386.4]
  wire [15:0] _T_54228; // @[Mux.scala 19:72:@26387.4]
  wire [15:0] _T_54243; // @[Mux.scala 19:72:@26402.4]
  wire [15:0] _T_54245; // @[Mux.scala 19:72:@26403.4]
  wire [15:0] _T_54260; // @[Mux.scala 19:72:@26418.4]
  wire [15:0] _T_54262; // @[Mux.scala 19:72:@26419.4]
  wire [15:0] _T_54277; // @[Mux.scala 19:72:@26434.4]
  wire [15:0] _T_54279; // @[Mux.scala 19:72:@26435.4]
  wire [15:0] _T_54294; // @[Mux.scala 19:72:@26450.4]
  wire [15:0] _T_54296; // @[Mux.scala 19:72:@26451.4]
  wire [15:0] _T_54311; // @[Mux.scala 19:72:@26466.4]
  wire [15:0] _T_54313; // @[Mux.scala 19:72:@26467.4]
  wire [15:0] _T_54314; // @[Mux.scala 19:72:@26468.4]
  wire [15:0] _T_54315; // @[Mux.scala 19:72:@26469.4]
  wire [15:0] _T_54316; // @[Mux.scala 19:72:@26470.4]
  wire [15:0] _T_54317; // @[Mux.scala 19:72:@26471.4]
  wire [15:0] _T_54318; // @[Mux.scala 19:72:@26472.4]
  wire [15:0] _T_54319; // @[Mux.scala 19:72:@26473.4]
  wire [15:0] _T_54320; // @[Mux.scala 19:72:@26474.4]
  wire [15:0] _T_54321; // @[Mux.scala 19:72:@26475.4]
  wire [15:0] _T_54322; // @[Mux.scala 19:72:@26476.4]
  wire [15:0] _T_54323; // @[Mux.scala 19:72:@26477.4]
  wire [15:0] _T_54324; // @[Mux.scala 19:72:@26478.4]
  wire [15:0] _T_54325; // @[Mux.scala 19:72:@26479.4]
  wire [15:0] _T_54326; // @[Mux.scala 19:72:@26480.4]
  wire [15:0] _T_54327; // @[Mux.scala 19:72:@26481.4]
  wire [15:0] _T_54328; // @[Mux.scala 19:72:@26482.4]
  wire [7:0] _T_54906; // @[Mux.scala 19:72:@26832.4]
  wire [7:0] _T_54913; // @[Mux.scala 19:72:@26839.4]
  wire [15:0] _T_54914; // @[Mux.scala 19:72:@26840.4]
  wire [15:0] _T_54916; // @[Mux.scala 19:72:@26841.4]
  wire [7:0] _T_54923; // @[Mux.scala 19:72:@26848.4]
  wire [7:0] _T_54930; // @[Mux.scala 19:72:@26855.4]
  wire [15:0] _T_54931; // @[Mux.scala 19:72:@26856.4]
  wire [15:0] _T_54933; // @[Mux.scala 19:72:@26857.4]
  wire [7:0] _T_54940; // @[Mux.scala 19:72:@26864.4]
  wire [7:0] _T_54947; // @[Mux.scala 19:72:@26871.4]
  wire [15:0] _T_54948; // @[Mux.scala 19:72:@26872.4]
  wire [15:0] _T_54950; // @[Mux.scala 19:72:@26873.4]
  wire [7:0] _T_54957; // @[Mux.scala 19:72:@26880.4]
  wire [7:0] _T_54964; // @[Mux.scala 19:72:@26887.4]
  wire [15:0] _T_54965; // @[Mux.scala 19:72:@26888.4]
  wire [15:0] _T_54967; // @[Mux.scala 19:72:@26889.4]
  wire [7:0] _T_54974; // @[Mux.scala 19:72:@26896.4]
  wire [7:0] _T_54981; // @[Mux.scala 19:72:@26903.4]
  wire [15:0] _T_54982; // @[Mux.scala 19:72:@26904.4]
  wire [15:0] _T_54984; // @[Mux.scala 19:72:@26905.4]
  wire [7:0] _T_54991; // @[Mux.scala 19:72:@26912.4]
  wire [7:0] _T_54998; // @[Mux.scala 19:72:@26919.4]
  wire [15:0] _T_54999; // @[Mux.scala 19:72:@26920.4]
  wire [15:0] _T_55001; // @[Mux.scala 19:72:@26921.4]
  wire [7:0] _T_55008; // @[Mux.scala 19:72:@26928.4]
  wire [7:0] _T_55015; // @[Mux.scala 19:72:@26935.4]
  wire [15:0] _T_55016; // @[Mux.scala 19:72:@26936.4]
  wire [15:0] _T_55018; // @[Mux.scala 19:72:@26937.4]
  wire [7:0] _T_55025; // @[Mux.scala 19:72:@26944.4]
  wire [7:0] _T_55032; // @[Mux.scala 19:72:@26951.4]
  wire [15:0] _T_55033; // @[Mux.scala 19:72:@26952.4]
  wire [15:0] _T_55035; // @[Mux.scala 19:72:@26953.4]
  wire [15:0] _T_55050; // @[Mux.scala 19:72:@26968.4]
  wire [15:0] _T_55052; // @[Mux.scala 19:72:@26969.4]
  wire [15:0] _T_55067; // @[Mux.scala 19:72:@26984.4]
  wire [15:0] _T_55069; // @[Mux.scala 19:72:@26985.4]
  wire [15:0] _T_55084; // @[Mux.scala 19:72:@27000.4]
  wire [15:0] _T_55086; // @[Mux.scala 19:72:@27001.4]
  wire [15:0] _T_55101; // @[Mux.scala 19:72:@27016.4]
  wire [15:0] _T_55103; // @[Mux.scala 19:72:@27017.4]
  wire [15:0] _T_55118; // @[Mux.scala 19:72:@27032.4]
  wire [15:0] _T_55120; // @[Mux.scala 19:72:@27033.4]
  wire [15:0] _T_55135; // @[Mux.scala 19:72:@27048.4]
  wire [15:0] _T_55137; // @[Mux.scala 19:72:@27049.4]
  wire [15:0] _T_55152; // @[Mux.scala 19:72:@27064.4]
  wire [15:0] _T_55154; // @[Mux.scala 19:72:@27065.4]
  wire [15:0] _T_55169; // @[Mux.scala 19:72:@27080.4]
  wire [15:0] _T_55171; // @[Mux.scala 19:72:@27081.4]
  wire [15:0] _T_55172; // @[Mux.scala 19:72:@27082.4]
  wire [15:0] _T_55173; // @[Mux.scala 19:72:@27083.4]
  wire [15:0] _T_55174; // @[Mux.scala 19:72:@27084.4]
  wire [15:0] _T_55175; // @[Mux.scala 19:72:@27085.4]
  wire [15:0] _T_55176; // @[Mux.scala 19:72:@27086.4]
  wire [15:0] _T_55177; // @[Mux.scala 19:72:@27087.4]
  wire [15:0] _T_55178; // @[Mux.scala 19:72:@27088.4]
  wire [15:0] _T_55179; // @[Mux.scala 19:72:@27089.4]
  wire [15:0] _T_55180; // @[Mux.scala 19:72:@27090.4]
  wire [15:0] _T_55181; // @[Mux.scala 19:72:@27091.4]
  wire [15:0] _T_55182; // @[Mux.scala 19:72:@27092.4]
  wire [15:0] _T_55183; // @[Mux.scala 19:72:@27093.4]
  wire [15:0] _T_55184; // @[Mux.scala 19:72:@27094.4]
  wire [15:0] _T_55185; // @[Mux.scala 19:72:@27095.4]
  wire [15:0] _T_55186; // @[Mux.scala 19:72:@27096.4]
  wire [7:0] _T_55764; // @[Mux.scala 19:72:@27446.4]
  wire [7:0] _T_55771; // @[Mux.scala 19:72:@27453.4]
  wire [15:0] _T_55772; // @[Mux.scala 19:72:@27454.4]
  wire [15:0] _T_55774; // @[Mux.scala 19:72:@27455.4]
  wire [7:0] _T_55781; // @[Mux.scala 19:72:@27462.4]
  wire [7:0] _T_55788; // @[Mux.scala 19:72:@27469.4]
  wire [15:0] _T_55789; // @[Mux.scala 19:72:@27470.4]
  wire [15:0] _T_55791; // @[Mux.scala 19:72:@27471.4]
  wire [7:0] _T_55798; // @[Mux.scala 19:72:@27478.4]
  wire [7:0] _T_55805; // @[Mux.scala 19:72:@27485.4]
  wire [15:0] _T_55806; // @[Mux.scala 19:72:@27486.4]
  wire [15:0] _T_55808; // @[Mux.scala 19:72:@27487.4]
  wire [7:0] _T_55815; // @[Mux.scala 19:72:@27494.4]
  wire [7:0] _T_55822; // @[Mux.scala 19:72:@27501.4]
  wire [15:0] _T_55823; // @[Mux.scala 19:72:@27502.4]
  wire [15:0] _T_55825; // @[Mux.scala 19:72:@27503.4]
  wire [7:0] _T_55832; // @[Mux.scala 19:72:@27510.4]
  wire [7:0] _T_55839; // @[Mux.scala 19:72:@27517.4]
  wire [15:0] _T_55840; // @[Mux.scala 19:72:@27518.4]
  wire [15:0] _T_55842; // @[Mux.scala 19:72:@27519.4]
  wire [7:0] _T_55849; // @[Mux.scala 19:72:@27526.4]
  wire [7:0] _T_55856; // @[Mux.scala 19:72:@27533.4]
  wire [15:0] _T_55857; // @[Mux.scala 19:72:@27534.4]
  wire [15:0] _T_55859; // @[Mux.scala 19:72:@27535.4]
  wire [7:0] _T_55866; // @[Mux.scala 19:72:@27542.4]
  wire [7:0] _T_55873; // @[Mux.scala 19:72:@27549.4]
  wire [15:0] _T_55874; // @[Mux.scala 19:72:@27550.4]
  wire [15:0] _T_55876; // @[Mux.scala 19:72:@27551.4]
  wire [7:0] _T_55883; // @[Mux.scala 19:72:@27558.4]
  wire [7:0] _T_55890; // @[Mux.scala 19:72:@27565.4]
  wire [15:0] _T_55891; // @[Mux.scala 19:72:@27566.4]
  wire [15:0] _T_55893; // @[Mux.scala 19:72:@27567.4]
  wire [15:0] _T_55908; // @[Mux.scala 19:72:@27582.4]
  wire [15:0] _T_55910; // @[Mux.scala 19:72:@27583.4]
  wire [15:0] _T_55925; // @[Mux.scala 19:72:@27598.4]
  wire [15:0] _T_55927; // @[Mux.scala 19:72:@27599.4]
  wire [15:0] _T_55942; // @[Mux.scala 19:72:@27614.4]
  wire [15:0] _T_55944; // @[Mux.scala 19:72:@27615.4]
  wire [15:0] _T_55959; // @[Mux.scala 19:72:@27630.4]
  wire [15:0] _T_55961; // @[Mux.scala 19:72:@27631.4]
  wire [15:0] _T_55976; // @[Mux.scala 19:72:@27646.4]
  wire [15:0] _T_55978; // @[Mux.scala 19:72:@27647.4]
  wire [15:0] _T_55993; // @[Mux.scala 19:72:@27662.4]
  wire [15:0] _T_55995; // @[Mux.scala 19:72:@27663.4]
  wire [15:0] _T_56010; // @[Mux.scala 19:72:@27678.4]
  wire [15:0] _T_56012; // @[Mux.scala 19:72:@27679.4]
  wire [15:0] _T_56027; // @[Mux.scala 19:72:@27694.4]
  wire [15:0] _T_56029; // @[Mux.scala 19:72:@27695.4]
  wire [15:0] _T_56030; // @[Mux.scala 19:72:@27696.4]
  wire [15:0] _T_56031; // @[Mux.scala 19:72:@27697.4]
  wire [15:0] _T_56032; // @[Mux.scala 19:72:@27698.4]
  wire [15:0] _T_56033; // @[Mux.scala 19:72:@27699.4]
  wire [15:0] _T_56034; // @[Mux.scala 19:72:@27700.4]
  wire [15:0] _T_56035; // @[Mux.scala 19:72:@27701.4]
  wire [15:0] _T_56036; // @[Mux.scala 19:72:@27702.4]
  wire [15:0] _T_56037; // @[Mux.scala 19:72:@27703.4]
  wire [15:0] _T_56038; // @[Mux.scala 19:72:@27704.4]
  wire [15:0] _T_56039; // @[Mux.scala 19:72:@27705.4]
  wire [15:0] _T_56040; // @[Mux.scala 19:72:@27706.4]
  wire [15:0] _T_56041; // @[Mux.scala 19:72:@27707.4]
  wire [15:0] _T_56042; // @[Mux.scala 19:72:@27708.4]
  wire [15:0] _T_56043; // @[Mux.scala 19:72:@27709.4]
  wire [15:0] _T_56044; // @[Mux.scala 19:72:@27710.4]
  wire [7:0] _T_56622; // @[Mux.scala 19:72:@28060.4]
  wire [7:0] _T_56629; // @[Mux.scala 19:72:@28067.4]
  wire [15:0] _T_56630; // @[Mux.scala 19:72:@28068.4]
  wire [15:0] _T_56632; // @[Mux.scala 19:72:@28069.4]
  wire [7:0] _T_56639; // @[Mux.scala 19:72:@28076.4]
  wire [7:0] _T_56646; // @[Mux.scala 19:72:@28083.4]
  wire [15:0] _T_56647; // @[Mux.scala 19:72:@28084.4]
  wire [15:0] _T_56649; // @[Mux.scala 19:72:@28085.4]
  wire [7:0] _T_56656; // @[Mux.scala 19:72:@28092.4]
  wire [7:0] _T_56663; // @[Mux.scala 19:72:@28099.4]
  wire [15:0] _T_56664; // @[Mux.scala 19:72:@28100.4]
  wire [15:0] _T_56666; // @[Mux.scala 19:72:@28101.4]
  wire [7:0] _T_56673; // @[Mux.scala 19:72:@28108.4]
  wire [7:0] _T_56680; // @[Mux.scala 19:72:@28115.4]
  wire [15:0] _T_56681; // @[Mux.scala 19:72:@28116.4]
  wire [15:0] _T_56683; // @[Mux.scala 19:72:@28117.4]
  wire [7:0] _T_56690; // @[Mux.scala 19:72:@28124.4]
  wire [7:0] _T_56697; // @[Mux.scala 19:72:@28131.4]
  wire [15:0] _T_56698; // @[Mux.scala 19:72:@28132.4]
  wire [15:0] _T_56700; // @[Mux.scala 19:72:@28133.4]
  wire [7:0] _T_56707; // @[Mux.scala 19:72:@28140.4]
  wire [7:0] _T_56714; // @[Mux.scala 19:72:@28147.4]
  wire [15:0] _T_56715; // @[Mux.scala 19:72:@28148.4]
  wire [15:0] _T_56717; // @[Mux.scala 19:72:@28149.4]
  wire [7:0] _T_56724; // @[Mux.scala 19:72:@28156.4]
  wire [7:0] _T_56731; // @[Mux.scala 19:72:@28163.4]
  wire [15:0] _T_56732; // @[Mux.scala 19:72:@28164.4]
  wire [15:0] _T_56734; // @[Mux.scala 19:72:@28165.4]
  wire [7:0] _T_56741; // @[Mux.scala 19:72:@28172.4]
  wire [7:0] _T_56748; // @[Mux.scala 19:72:@28179.4]
  wire [15:0] _T_56749; // @[Mux.scala 19:72:@28180.4]
  wire [15:0] _T_56751; // @[Mux.scala 19:72:@28181.4]
  wire [15:0] _T_56766; // @[Mux.scala 19:72:@28196.4]
  wire [15:0] _T_56768; // @[Mux.scala 19:72:@28197.4]
  wire [15:0] _T_56783; // @[Mux.scala 19:72:@28212.4]
  wire [15:0] _T_56785; // @[Mux.scala 19:72:@28213.4]
  wire [15:0] _T_56800; // @[Mux.scala 19:72:@28228.4]
  wire [15:0] _T_56802; // @[Mux.scala 19:72:@28229.4]
  wire [15:0] _T_56817; // @[Mux.scala 19:72:@28244.4]
  wire [15:0] _T_56819; // @[Mux.scala 19:72:@28245.4]
  wire [15:0] _T_56834; // @[Mux.scala 19:72:@28260.4]
  wire [15:0] _T_56836; // @[Mux.scala 19:72:@28261.4]
  wire [15:0] _T_56851; // @[Mux.scala 19:72:@28276.4]
  wire [15:0] _T_56853; // @[Mux.scala 19:72:@28277.4]
  wire [15:0] _T_56868; // @[Mux.scala 19:72:@28292.4]
  wire [15:0] _T_56870; // @[Mux.scala 19:72:@28293.4]
  wire [15:0] _T_56885; // @[Mux.scala 19:72:@28308.4]
  wire [15:0] _T_56887; // @[Mux.scala 19:72:@28309.4]
  wire [15:0] _T_56888; // @[Mux.scala 19:72:@28310.4]
  wire [15:0] _T_56889; // @[Mux.scala 19:72:@28311.4]
  wire [15:0] _T_56890; // @[Mux.scala 19:72:@28312.4]
  wire [15:0] _T_56891; // @[Mux.scala 19:72:@28313.4]
  wire [15:0] _T_56892; // @[Mux.scala 19:72:@28314.4]
  wire [15:0] _T_56893; // @[Mux.scala 19:72:@28315.4]
  wire [15:0] _T_56894; // @[Mux.scala 19:72:@28316.4]
  wire [15:0] _T_56895; // @[Mux.scala 19:72:@28317.4]
  wire [15:0] _T_56896; // @[Mux.scala 19:72:@28318.4]
  wire [15:0] _T_56897; // @[Mux.scala 19:72:@28319.4]
  wire [15:0] _T_56898; // @[Mux.scala 19:72:@28320.4]
  wire [15:0] _T_56899; // @[Mux.scala 19:72:@28321.4]
  wire [15:0] _T_56900; // @[Mux.scala 19:72:@28322.4]
  wire [15:0] _T_56901; // @[Mux.scala 19:72:@28323.4]
  wire [15:0] _T_56902; // @[Mux.scala 19:72:@28324.4]
  wire [7:0] _T_57480; // @[Mux.scala 19:72:@28674.4]
  wire [7:0] _T_57487; // @[Mux.scala 19:72:@28681.4]
  wire [15:0] _T_57488; // @[Mux.scala 19:72:@28682.4]
  wire [15:0] _T_57490; // @[Mux.scala 19:72:@28683.4]
  wire [7:0] _T_57497; // @[Mux.scala 19:72:@28690.4]
  wire [7:0] _T_57504; // @[Mux.scala 19:72:@28697.4]
  wire [15:0] _T_57505; // @[Mux.scala 19:72:@28698.4]
  wire [15:0] _T_57507; // @[Mux.scala 19:72:@28699.4]
  wire [7:0] _T_57514; // @[Mux.scala 19:72:@28706.4]
  wire [7:0] _T_57521; // @[Mux.scala 19:72:@28713.4]
  wire [15:0] _T_57522; // @[Mux.scala 19:72:@28714.4]
  wire [15:0] _T_57524; // @[Mux.scala 19:72:@28715.4]
  wire [7:0] _T_57531; // @[Mux.scala 19:72:@28722.4]
  wire [7:0] _T_57538; // @[Mux.scala 19:72:@28729.4]
  wire [15:0] _T_57539; // @[Mux.scala 19:72:@28730.4]
  wire [15:0] _T_57541; // @[Mux.scala 19:72:@28731.4]
  wire [7:0] _T_57548; // @[Mux.scala 19:72:@28738.4]
  wire [7:0] _T_57555; // @[Mux.scala 19:72:@28745.4]
  wire [15:0] _T_57556; // @[Mux.scala 19:72:@28746.4]
  wire [15:0] _T_57558; // @[Mux.scala 19:72:@28747.4]
  wire [7:0] _T_57565; // @[Mux.scala 19:72:@28754.4]
  wire [7:0] _T_57572; // @[Mux.scala 19:72:@28761.4]
  wire [15:0] _T_57573; // @[Mux.scala 19:72:@28762.4]
  wire [15:0] _T_57575; // @[Mux.scala 19:72:@28763.4]
  wire [7:0] _T_57582; // @[Mux.scala 19:72:@28770.4]
  wire [7:0] _T_57589; // @[Mux.scala 19:72:@28777.4]
  wire [15:0] _T_57590; // @[Mux.scala 19:72:@28778.4]
  wire [15:0] _T_57592; // @[Mux.scala 19:72:@28779.4]
  wire [7:0] _T_57599; // @[Mux.scala 19:72:@28786.4]
  wire [7:0] _T_57606; // @[Mux.scala 19:72:@28793.4]
  wire [15:0] _T_57607; // @[Mux.scala 19:72:@28794.4]
  wire [15:0] _T_57609; // @[Mux.scala 19:72:@28795.4]
  wire [15:0] _T_57624; // @[Mux.scala 19:72:@28810.4]
  wire [15:0] _T_57626; // @[Mux.scala 19:72:@28811.4]
  wire [15:0] _T_57641; // @[Mux.scala 19:72:@28826.4]
  wire [15:0] _T_57643; // @[Mux.scala 19:72:@28827.4]
  wire [15:0] _T_57658; // @[Mux.scala 19:72:@28842.4]
  wire [15:0] _T_57660; // @[Mux.scala 19:72:@28843.4]
  wire [15:0] _T_57675; // @[Mux.scala 19:72:@28858.4]
  wire [15:0] _T_57677; // @[Mux.scala 19:72:@28859.4]
  wire [15:0] _T_57692; // @[Mux.scala 19:72:@28874.4]
  wire [15:0] _T_57694; // @[Mux.scala 19:72:@28875.4]
  wire [15:0] _T_57709; // @[Mux.scala 19:72:@28890.4]
  wire [15:0] _T_57711; // @[Mux.scala 19:72:@28891.4]
  wire [15:0] _T_57726; // @[Mux.scala 19:72:@28906.4]
  wire [15:0] _T_57728; // @[Mux.scala 19:72:@28907.4]
  wire [15:0] _T_57743; // @[Mux.scala 19:72:@28922.4]
  wire [15:0] _T_57745; // @[Mux.scala 19:72:@28923.4]
  wire [15:0] _T_57746; // @[Mux.scala 19:72:@28924.4]
  wire [15:0] _T_57747; // @[Mux.scala 19:72:@28925.4]
  wire [15:0] _T_57748; // @[Mux.scala 19:72:@28926.4]
  wire [15:0] _T_57749; // @[Mux.scala 19:72:@28927.4]
  wire [15:0] _T_57750; // @[Mux.scala 19:72:@28928.4]
  wire [15:0] _T_57751; // @[Mux.scala 19:72:@28929.4]
  wire [15:0] _T_57752; // @[Mux.scala 19:72:@28930.4]
  wire [15:0] _T_57753; // @[Mux.scala 19:72:@28931.4]
  wire [15:0] _T_57754; // @[Mux.scala 19:72:@28932.4]
  wire [15:0] _T_57755; // @[Mux.scala 19:72:@28933.4]
  wire [15:0] _T_57756; // @[Mux.scala 19:72:@28934.4]
  wire [15:0] _T_57757; // @[Mux.scala 19:72:@28935.4]
  wire [15:0] _T_57758; // @[Mux.scala 19:72:@28936.4]
  wire [15:0] _T_57759; // @[Mux.scala 19:72:@28937.4]
  wire [15:0] _T_57760; // @[Mux.scala 19:72:@28938.4]
  wire [7:0] _T_58338; // @[Mux.scala 19:72:@29288.4]
  wire [7:0] _T_58345; // @[Mux.scala 19:72:@29295.4]
  wire [15:0] _T_58346; // @[Mux.scala 19:72:@29296.4]
  wire [15:0] _T_58348; // @[Mux.scala 19:72:@29297.4]
  wire [7:0] _T_58355; // @[Mux.scala 19:72:@29304.4]
  wire [7:0] _T_58362; // @[Mux.scala 19:72:@29311.4]
  wire [15:0] _T_58363; // @[Mux.scala 19:72:@29312.4]
  wire [15:0] _T_58365; // @[Mux.scala 19:72:@29313.4]
  wire [7:0] _T_58372; // @[Mux.scala 19:72:@29320.4]
  wire [7:0] _T_58379; // @[Mux.scala 19:72:@29327.4]
  wire [15:0] _T_58380; // @[Mux.scala 19:72:@29328.4]
  wire [15:0] _T_58382; // @[Mux.scala 19:72:@29329.4]
  wire [7:0] _T_58389; // @[Mux.scala 19:72:@29336.4]
  wire [7:0] _T_58396; // @[Mux.scala 19:72:@29343.4]
  wire [15:0] _T_58397; // @[Mux.scala 19:72:@29344.4]
  wire [15:0] _T_58399; // @[Mux.scala 19:72:@29345.4]
  wire [7:0] _T_58406; // @[Mux.scala 19:72:@29352.4]
  wire [7:0] _T_58413; // @[Mux.scala 19:72:@29359.4]
  wire [15:0] _T_58414; // @[Mux.scala 19:72:@29360.4]
  wire [15:0] _T_58416; // @[Mux.scala 19:72:@29361.4]
  wire [7:0] _T_58423; // @[Mux.scala 19:72:@29368.4]
  wire [7:0] _T_58430; // @[Mux.scala 19:72:@29375.4]
  wire [15:0] _T_58431; // @[Mux.scala 19:72:@29376.4]
  wire [15:0] _T_58433; // @[Mux.scala 19:72:@29377.4]
  wire [7:0] _T_58440; // @[Mux.scala 19:72:@29384.4]
  wire [7:0] _T_58447; // @[Mux.scala 19:72:@29391.4]
  wire [15:0] _T_58448; // @[Mux.scala 19:72:@29392.4]
  wire [15:0] _T_58450; // @[Mux.scala 19:72:@29393.4]
  wire [7:0] _T_58457; // @[Mux.scala 19:72:@29400.4]
  wire [7:0] _T_58464; // @[Mux.scala 19:72:@29407.4]
  wire [15:0] _T_58465; // @[Mux.scala 19:72:@29408.4]
  wire [15:0] _T_58467; // @[Mux.scala 19:72:@29409.4]
  wire [15:0] _T_58482; // @[Mux.scala 19:72:@29424.4]
  wire [15:0] _T_58484; // @[Mux.scala 19:72:@29425.4]
  wire [15:0] _T_58499; // @[Mux.scala 19:72:@29440.4]
  wire [15:0] _T_58501; // @[Mux.scala 19:72:@29441.4]
  wire [15:0] _T_58516; // @[Mux.scala 19:72:@29456.4]
  wire [15:0] _T_58518; // @[Mux.scala 19:72:@29457.4]
  wire [15:0] _T_58533; // @[Mux.scala 19:72:@29472.4]
  wire [15:0] _T_58535; // @[Mux.scala 19:72:@29473.4]
  wire [15:0] _T_58550; // @[Mux.scala 19:72:@29488.4]
  wire [15:0] _T_58552; // @[Mux.scala 19:72:@29489.4]
  wire [15:0] _T_58567; // @[Mux.scala 19:72:@29504.4]
  wire [15:0] _T_58569; // @[Mux.scala 19:72:@29505.4]
  wire [15:0] _T_58584; // @[Mux.scala 19:72:@29520.4]
  wire [15:0] _T_58586; // @[Mux.scala 19:72:@29521.4]
  wire [15:0] _T_58601; // @[Mux.scala 19:72:@29536.4]
  wire [15:0] _T_58603; // @[Mux.scala 19:72:@29537.4]
  wire [15:0] _T_58604; // @[Mux.scala 19:72:@29538.4]
  wire [15:0] _T_58605; // @[Mux.scala 19:72:@29539.4]
  wire [15:0] _T_58606; // @[Mux.scala 19:72:@29540.4]
  wire [15:0] _T_58607; // @[Mux.scala 19:72:@29541.4]
  wire [15:0] _T_58608; // @[Mux.scala 19:72:@29542.4]
  wire [15:0] _T_58609; // @[Mux.scala 19:72:@29543.4]
  wire [15:0] _T_58610; // @[Mux.scala 19:72:@29544.4]
  wire [15:0] _T_58611; // @[Mux.scala 19:72:@29545.4]
  wire [15:0] _T_58612; // @[Mux.scala 19:72:@29546.4]
  wire [15:0] _T_58613; // @[Mux.scala 19:72:@29547.4]
  wire [15:0] _T_58614; // @[Mux.scala 19:72:@29548.4]
  wire [15:0] _T_58615; // @[Mux.scala 19:72:@29549.4]
  wire [15:0] _T_58616; // @[Mux.scala 19:72:@29550.4]
  wire [15:0] _T_58617; // @[Mux.scala 19:72:@29551.4]
  wire [15:0] _T_58618; // @[Mux.scala 19:72:@29552.4]
  wire [7:0] _T_59196; // @[Mux.scala 19:72:@29902.4]
  wire [7:0] _T_59203; // @[Mux.scala 19:72:@29909.4]
  wire [15:0] _T_59204; // @[Mux.scala 19:72:@29910.4]
  wire [15:0] _T_59206; // @[Mux.scala 19:72:@29911.4]
  wire [7:0] _T_59213; // @[Mux.scala 19:72:@29918.4]
  wire [7:0] _T_59220; // @[Mux.scala 19:72:@29925.4]
  wire [15:0] _T_59221; // @[Mux.scala 19:72:@29926.4]
  wire [15:0] _T_59223; // @[Mux.scala 19:72:@29927.4]
  wire [7:0] _T_59230; // @[Mux.scala 19:72:@29934.4]
  wire [7:0] _T_59237; // @[Mux.scala 19:72:@29941.4]
  wire [15:0] _T_59238; // @[Mux.scala 19:72:@29942.4]
  wire [15:0] _T_59240; // @[Mux.scala 19:72:@29943.4]
  wire [7:0] _T_59247; // @[Mux.scala 19:72:@29950.4]
  wire [7:0] _T_59254; // @[Mux.scala 19:72:@29957.4]
  wire [15:0] _T_59255; // @[Mux.scala 19:72:@29958.4]
  wire [15:0] _T_59257; // @[Mux.scala 19:72:@29959.4]
  wire [7:0] _T_59264; // @[Mux.scala 19:72:@29966.4]
  wire [7:0] _T_59271; // @[Mux.scala 19:72:@29973.4]
  wire [15:0] _T_59272; // @[Mux.scala 19:72:@29974.4]
  wire [15:0] _T_59274; // @[Mux.scala 19:72:@29975.4]
  wire [7:0] _T_59281; // @[Mux.scala 19:72:@29982.4]
  wire [7:0] _T_59288; // @[Mux.scala 19:72:@29989.4]
  wire [15:0] _T_59289; // @[Mux.scala 19:72:@29990.4]
  wire [15:0] _T_59291; // @[Mux.scala 19:72:@29991.4]
  wire [7:0] _T_59298; // @[Mux.scala 19:72:@29998.4]
  wire [7:0] _T_59305; // @[Mux.scala 19:72:@30005.4]
  wire [15:0] _T_59306; // @[Mux.scala 19:72:@30006.4]
  wire [15:0] _T_59308; // @[Mux.scala 19:72:@30007.4]
  wire [7:0] _T_59315; // @[Mux.scala 19:72:@30014.4]
  wire [7:0] _T_59322; // @[Mux.scala 19:72:@30021.4]
  wire [15:0] _T_59323; // @[Mux.scala 19:72:@30022.4]
  wire [15:0] _T_59325; // @[Mux.scala 19:72:@30023.4]
  wire [15:0] _T_59340; // @[Mux.scala 19:72:@30038.4]
  wire [15:0] _T_59342; // @[Mux.scala 19:72:@30039.4]
  wire [15:0] _T_59357; // @[Mux.scala 19:72:@30054.4]
  wire [15:0] _T_59359; // @[Mux.scala 19:72:@30055.4]
  wire [15:0] _T_59374; // @[Mux.scala 19:72:@30070.4]
  wire [15:0] _T_59376; // @[Mux.scala 19:72:@30071.4]
  wire [15:0] _T_59391; // @[Mux.scala 19:72:@30086.4]
  wire [15:0] _T_59393; // @[Mux.scala 19:72:@30087.4]
  wire [15:0] _T_59408; // @[Mux.scala 19:72:@30102.4]
  wire [15:0] _T_59410; // @[Mux.scala 19:72:@30103.4]
  wire [15:0] _T_59425; // @[Mux.scala 19:72:@30118.4]
  wire [15:0] _T_59427; // @[Mux.scala 19:72:@30119.4]
  wire [15:0] _T_59442; // @[Mux.scala 19:72:@30134.4]
  wire [15:0] _T_59444; // @[Mux.scala 19:72:@30135.4]
  wire [15:0] _T_59459; // @[Mux.scala 19:72:@30150.4]
  wire [15:0] _T_59461; // @[Mux.scala 19:72:@30151.4]
  wire [15:0] _T_59462; // @[Mux.scala 19:72:@30152.4]
  wire [15:0] _T_59463; // @[Mux.scala 19:72:@30153.4]
  wire [15:0] _T_59464; // @[Mux.scala 19:72:@30154.4]
  wire [15:0] _T_59465; // @[Mux.scala 19:72:@30155.4]
  wire [15:0] _T_59466; // @[Mux.scala 19:72:@30156.4]
  wire [15:0] _T_59467; // @[Mux.scala 19:72:@30157.4]
  wire [15:0] _T_59468; // @[Mux.scala 19:72:@30158.4]
  wire [15:0] _T_59469; // @[Mux.scala 19:72:@30159.4]
  wire [15:0] _T_59470; // @[Mux.scala 19:72:@30160.4]
  wire [15:0] _T_59471; // @[Mux.scala 19:72:@30161.4]
  wire [15:0] _T_59472; // @[Mux.scala 19:72:@30162.4]
  wire [15:0] _T_59473; // @[Mux.scala 19:72:@30163.4]
  wire [15:0] _T_59474; // @[Mux.scala 19:72:@30164.4]
  wire [15:0] _T_59475; // @[Mux.scala 19:72:@30165.4]
  wire [15:0] _T_59476; // @[Mux.scala 19:72:@30166.4]
  wire [7:0] _T_60054; // @[Mux.scala 19:72:@30516.4]
  wire [7:0] _T_60061; // @[Mux.scala 19:72:@30523.4]
  wire [15:0] _T_60062; // @[Mux.scala 19:72:@30524.4]
  wire [15:0] _T_60064; // @[Mux.scala 19:72:@30525.4]
  wire [7:0] _T_60071; // @[Mux.scala 19:72:@30532.4]
  wire [7:0] _T_60078; // @[Mux.scala 19:72:@30539.4]
  wire [15:0] _T_60079; // @[Mux.scala 19:72:@30540.4]
  wire [15:0] _T_60081; // @[Mux.scala 19:72:@30541.4]
  wire [7:0] _T_60088; // @[Mux.scala 19:72:@30548.4]
  wire [7:0] _T_60095; // @[Mux.scala 19:72:@30555.4]
  wire [15:0] _T_60096; // @[Mux.scala 19:72:@30556.4]
  wire [15:0] _T_60098; // @[Mux.scala 19:72:@30557.4]
  wire [7:0] _T_60105; // @[Mux.scala 19:72:@30564.4]
  wire [7:0] _T_60112; // @[Mux.scala 19:72:@30571.4]
  wire [15:0] _T_60113; // @[Mux.scala 19:72:@30572.4]
  wire [15:0] _T_60115; // @[Mux.scala 19:72:@30573.4]
  wire [7:0] _T_60122; // @[Mux.scala 19:72:@30580.4]
  wire [7:0] _T_60129; // @[Mux.scala 19:72:@30587.4]
  wire [15:0] _T_60130; // @[Mux.scala 19:72:@30588.4]
  wire [15:0] _T_60132; // @[Mux.scala 19:72:@30589.4]
  wire [7:0] _T_60139; // @[Mux.scala 19:72:@30596.4]
  wire [7:0] _T_60146; // @[Mux.scala 19:72:@30603.4]
  wire [15:0] _T_60147; // @[Mux.scala 19:72:@30604.4]
  wire [15:0] _T_60149; // @[Mux.scala 19:72:@30605.4]
  wire [7:0] _T_60156; // @[Mux.scala 19:72:@30612.4]
  wire [7:0] _T_60163; // @[Mux.scala 19:72:@30619.4]
  wire [15:0] _T_60164; // @[Mux.scala 19:72:@30620.4]
  wire [15:0] _T_60166; // @[Mux.scala 19:72:@30621.4]
  wire [7:0] _T_60173; // @[Mux.scala 19:72:@30628.4]
  wire [7:0] _T_60180; // @[Mux.scala 19:72:@30635.4]
  wire [15:0] _T_60181; // @[Mux.scala 19:72:@30636.4]
  wire [15:0] _T_60183; // @[Mux.scala 19:72:@30637.4]
  wire [15:0] _T_60198; // @[Mux.scala 19:72:@30652.4]
  wire [15:0] _T_60200; // @[Mux.scala 19:72:@30653.4]
  wire [15:0] _T_60215; // @[Mux.scala 19:72:@30668.4]
  wire [15:0] _T_60217; // @[Mux.scala 19:72:@30669.4]
  wire [15:0] _T_60232; // @[Mux.scala 19:72:@30684.4]
  wire [15:0] _T_60234; // @[Mux.scala 19:72:@30685.4]
  wire [15:0] _T_60249; // @[Mux.scala 19:72:@30700.4]
  wire [15:0] _T_60251; // @[Mux.scala 19:72:@30701.4]
  wire [15:0] _T_60266; // @[Mux.scala 19:72:@30716.4]
  wire [15:0] _T_60268; // @[Mux.scala 19:72:@30717.4]
  wire [15:0] _T_60283; // @[Mux.scala 19:72:@30732.4]
  wire [15:0] _T_60285; // @[Mux.scala 19:72:@30733.4]
  wire [15:0] _T_60300; // @[Mux.scala 19:72:@30748.4]
  wire [15:0] _T_60302; // @[Mux.scala 19:72:@30749.4]
  wire [15:0] _T_60317; // @[Mux.scala 19:72:@30764.4]
  wire [15:0] _T_60319; // @[Mux.scala 19:72:@30765.4]
  wire [15:0] _T_60320; // @[Mux.scala 19:72:@30766.4]
  wire [15:0] _T_60321; // @[Mux.scala 19:72:@30767.4]
  wire [15:0] _T_60322; // @[Mux.scala 19:72:@30768.4]
  wire [15:0] _T_60323; // @[Mux.scala 19:72:@30769.4]
  wire [15:0] _T_60324; // @[Mux.scala 19:72:@30770.4]
  wire [15:0] _T_60325; // @[Mux.scala 19:72:@30771.4]
  wire [15:0] _T_60326; // @[Mux.scala 19:72:@30772.4]
  wire [15:0] _T_60327; // @[Mux.scala 19:72:@30773.4]
  wire [15:0] _T_60328; // @[Mux.scala 19:72:@30774.4]
  wire [15:0] _T_60329; // @[Mux.scala 19:72:@30775.4]
  wire [15:0] _T_60330; // @[Mux.scala 19:72:@30776.4]
  wire [15:0] _T_60331; // @[Mux.scala 19:72:@30777.4]
  wire [15:0] _T_60332; // @[Mux.scala 19:72:@30778.4]
  wire [15:0] _T_60333; // @[Mux.scala 19:72:@30779.4]
  wire [15:0] _T_60334; // @[Mux.scala 19:72:@30780.4]
  wire [7:0] _T_60912; // @[Mux.scala 19:72:@31130.4]
  wire [7:0] _T_60919; // @[Mux.scala 19:72:@31137.4]
  wire [15:0] _T_60920; // @[Mux.scala 19:72:@31138.4]
  wire [15:0] _T_60922; // @[Mux.scala 19:72:@31139.4]
  wire [7:0] _T_60929; // @[Mux.scala 19:72:@31146.4]
  wire [7:0] _T_60936; // @[Mux.scala 19:72:@31153.4]
  wire [15:0] _T_60937; // @[Mux.scala 19:72:@31154.4]
  wire [15:0] _T_60939; // @[Mux.scala 19:72:@31155.4]
  wire [7:0] _T_60946; // @[Mux.scala 19:72:@31162.4]
  wire [7:0] _T_60953; // @[Mux.scala 19:72:@31169.4]
  wire [15:0] _T_60954; // @[Mux.scala 19:72:@31170.4]
  wire [15:0] _T_60956; // @[Mux.scala 19:72:@31171.4]
  wire [7:0] _T_60963; // @[Mux.scala 19:72:@31178.4]
  wire [7:0] _T_60970; // @[Mux.scala 19:72:@31185.4]
  wire [15:0] _T_60971; // @[Mux.scala 19:72:@31186.4]
  wire [15:0] _T_60973; // @[Mux.scala 19:72:@31187.4]
  wire [7:0] _T_60980; // @[Mux.scala 19:72:@31194.4]
  wire [7:0] _T_60987; // @[Mux.scala 19:72:@31201.4]
  wire [15:0] _T_60988; // @[Mux.scala 19:72:@31202.4]
  wire [15:0] _T_60990; // @[Mux.scala 19:72:@31203.4]
  wire [7:0] _T_60997; // @[Mux.scala 19:72:@31210.4]
  wire [7:0] _T_61004; // @[Mux.scala 19:72:@31217.4]
  wire [15:0] _T_61005; // @[Mux.scala 19:72:@31218.4]
  wire [15:0] _T_61007; // @[Mux.scala 19:72:@31219.4]
  wire [7:0] _T_61014; // @[Mux.scala 19:72:@31226.4]
  wire [7:0] _T_61021; // @[Mux.scala 19:72:@31233.4]
  wire [15:0] _T_61022; // @[Mux.scala 19:72:@31234.4]
  wire [15:0] _T_61024; // @[Mux.scala 19:72:@31235.4]
  wire [7:0] _T_61031; // @[Mux.scala 19:72:@31242.4]
  wire [7:0] _T_61038; // @[Mux.scala 19:72:@31249.4]
  wire [15:0] _T_61039; // @[Mux.scala 19:72:@31250.4]
  wire [15:0] _T_61041; // @[Mux.scala 19:72:@31251.4]
  wire [15:0] _T_61056; // @[Mux.scala 19:72:@31266.4]
  wire [15:0] _T_61058; // @[Mux.scala 19:72:@31267.4]
  wire [15:0] _T_61073; // @[Mux.scala 19:72:@31282.4]
  wire [15:0] _T_61075; // @[Mux.scala 19:72:@31283.4]
  wire [15:0] _T_61090; // @[Mux.scala 19:72:@31298.4]
  wire [15:0] _T_61092; // @[Mux.scala 19:72:@31299.4]
  wire [15:0] _T_61107; // @[Mux.scala 19:72:@31314.4]
  wire [15:0] _T_61109; // @[Mux.scala 19:72:@31315.4]
  wire [15:0] _T_61124; // @[Mux.scala 19:72:@31330.4]
  wire [15:0] _T_61126; // @[Mux.scala 19:72:@31331.4]
  wire [15:0] _T_61141; // @[Mux.scala 19:72:@31346.4]
  wire [15:0] _T_61143; // @[Mux.scala 19:72:@31347.4]
  wire [15:0] _T_61158; // @[Mux.scala 19:72:@31362.4]
  wire [15:0] _T_61160; // @[Mux.scala 19:72:@31363.4]
  wire [15:0] _T_61175; // @[Mux.scala 19:72:@31378.4]
  wire [15:0] _T_61177; // @[Mux.scala 19:72:@31379.4]
  wire [15:0] _T_61178; // @[Mux.scala 19:72:@31380.4]
  wire [15:0] _T_61179; // @[Mux.scala 19:72:@31381.4]
  wire [15:0] _T_61180; // @[Mux.scala 19:72:@31382.4]
  wire [15:0] _T_61181; // @[Mux.scala 19:72:@31383.4]
  wire [15:0] _T_61182; // @[Mux.scala 19:72:@31384.4]
  wire [15:0] _T_61183; // @[Mux.scala 19:72:@31385.4]
  wire [15:0] _T_61184; // @[Mux.scala 19:72:@31386.4]
  wire [15:0] _T_61185; // @[Mux.scala 19:72:@31387.4]
  wire [15:0] _T_61186; // @[Mux.scala 19:72:@31388.4]
  wire [15:0] _T_61187; // @[Mux.scala 19:72:@31389.4]
  wire [15:0] _T_61188; // @[Mux.scala 19:72:@31390.4]
  wire [15:0] _T_61189; // @[Mux.scala 19:72:@31391.4]
  wire [15:0] _T_61190; // @[Mux.scala 19:72:@31392.4]
  wire [15:0] _T_61191; // @[Mux.scala 19:72:@31393.4]
  wire [15:0] _T_61192; // @[Mux.scala 19:72:@31394.4]
  wire [7:0] _T_61770; // @[Mux.scala 19:72:@31744.4]
  wire [7:0] _T_61777; // @[Mux.scala 19:72:@31751.4]
  wire [15:0] _T_61778; // @[Mux.scala 19:72:@31752.4]
  wire [15:0] _T_61780; // @[Mux.scala 19:72:@31753.4]
  wire [7:0] _T_61787; // @[Mux.scala 19:72:@31760.4]
  wire [7:0] _T_61794; // @[Mux.scala 19:72:@31767.4]
  wire [15:0] _T_61795; // @[Mux.scala 19:72:@31768.4]
  wire [15:0] _T_61797; // @[Mux.scala 19:72:@31769.4]
  wire [7:0] _T_61804; // @[Mux.scala 19:72:@31776.4]
  wire [7:0] _T_61811; // @[Mux.scala 19:72:@31783.4]
  wire [15:0] _T_61812; // @[Mux.scala 19:72:@31784.4]
  wire [15:0] _T_61814; // @[Mux.scala 19:72:@31785.4]
  wire [7:0] _T_61821; // @[Mux.scala 19:72:@31792.4]
  wire [7:0] _T_61828; // @[Mux.scala 19:72:@31799.4]
  wire [15:0] _T_61829; // @[Mux.scala 19:72:@31800.4]
  wire [15:0] _T_61831; // @[Mux.scala 19:72:@31801.4]
  wire [7:0] _T_61838; // @[Mux.scala 19:72:@31808.4]
  wire [7:0] _T_61845; // @[Mux.scala 19:72:@31815.4]
  wire [15:0] _T_61846; // @[Mux.scala 19:72:@31816.4]
  wire [15:0] _T_61848; // @[Mux.scala 19:72:@31817.4]
  wire [7:0] _T_61855; // @[Mux.scala 19:72:@31824.4]
  wire [7:0] _T_61862; // @[Mux.scala 19:72:@31831.4]
  wire [15:0] _T_61863; // @[Mux.scala 19:72:@31832.4]
  wire [15:0] _T_61865; // @[Mux.scala 19:72:@31833.4]
  wire [7:0] _T_61872; // @[Mux.scala 19:72:@31840.4]
  wire [7:0] _T_61879; // @[Mux.scala 19:72:@31847.4]
  wire [15:0] _T_61880; // @[Mux.scala 19:72:@31848.4]
  wire [15:0] _T_61882; // @[Mux.scala 19:72:@31849.4]
  wire [7:0] _T_61889; // @[Mux.scala 19:72:@31856.4]
  wire [7:0] _T_61896; // @[Mux.scala 19:72:@31863.4]
  wire [15:0] _T_61897; // @[Mux.scala 19:72:@31864.4]
  wire [15:0] _T_61899; // @[Mux.scala 19:72:@31865.4]
  wire [15:0] _T_61914; // @[Mux.scala 19:72:@31880.4]
  wire [15:0] _T_61916; // @[Mux.scala 19:72:@31881.4]
  wire [15:0] _T_61931; // @[Mux.scala 19:72:@31896.4]
  wire [15:0] _T_61933; // @[Mux.scala 19:72:@31897.4]
  wire [15:0] _T_61948; // @[Mux.scala 19:72:@31912.4]
  wire [15:0] _T_61950; // @[Mux.scala 19:72:@31913.4]
  wire [15:0] _T_61965; // @[Mux.scala 19:72:@31928.4]
  wire [15:0] _T_61967; // @[Mux.scala 19:72:@31929.4]
  wire [15:0] _T_61982; // @[Mux.scala 19:72:@31944.4]
  wire [15:0] _T_61984; // @[Mux.scala 19:72:@31945.4]
  wire [15:0] _T_61999; // @[Mux.scala 19:72:@31960.4]
  wire [15:0] _T_62001; // @[Mux.scala 19:72:@31961.4]
  wire [15:0] _T_62016; // @[Mux.scala 19:72:@31976.4]
  wire [15:0] _T_62018; // @[Mux.scala 19:72:@31977.4]
  wire [15:0] _T_62033; // @[Mux.scala 19:72:@31992.4]
  wire [15:0] _T_62035; // @[Mux.scala 19:72:@31993.4]
  wire [15:0] _T_62036; // @[Mux.scala 19:72:@31994.4]
  wire [15:0] _T_62037; // @[Mux.scala 19:72:@31995.4]
  wire [15:0] _T_62038; // @[Mux.scala 19:72:@31996.4]
  wire [15:0] _T_62039; // @[Mux.scala 19:72:@31997.4]
  wire [15:0] _T_62040; // @[Mux.scala 19:72:@31998.4]
  wire [15:0] _T_62041; // @[Mux.scala 19:72:@31999.4]
  wire [15:0] _T_62042; // @[Mux.scala 19:72:@32000.4]
  wire [15:0] _T_62043; // @[Mux.scala 19:72:@32001.4]
  wire [15:0] _T_62044; // @[Mux.scala 19:72:@32002.4]
  wire [15:0] _T_62045; // @[Mux.scala 19:72:@32003.4]
  wire [15:0] _T_62046; // @[Mux.scala 19:72:@32004.4]
  wire [15:0] _T_62047; // @[Mux.scala 19:72:@32005.4]
  wire [15:0] _T_62048; // @[Mux.scala 19:72:@32006.4]
  wire [15:0] _T_62049; // @[Mux.scala 19:72:@32007.4]
  wire [15:0] _T_62050; // @[Mux.scala 19:72:@32008.4]
  wire [7:0] _T_62628; // @[Mux.scala 19:72:@32358.4]
  wire [7:0] _T_62635; // @[Mux.scala 19:72:@32365.4]
  wire [15:0] _T_62636; // @[Mux.scala 19:72:@32366.4]
  wire [15:0] _T_62638; // @[Mux.scala 19:72:@32367.4]
  wire [7:0] _T_62645; // @[Mux.scala 19:72:@32374.4]
  wire [7:0] _T_62652; // @[Mux.scala 19:72:@32381.4]
  wire [15:0] _T_62653; // @[Mux.scala 19:72:@32382.4]
  wire [15:0] _T_62655; // @[Mux.scala 19:72:@32383.4]
  wire [7:0] _T_62662; // @[Mux.scala 19:72:@32390.4]
  wire [7:0] _T_62669; // @[Mux.scala 19:72:@32397.4]
  wire [15:0] _T_62670; // @[Mux.scala 19:72:@32398.4]
  wire [15:0] _T_62672; // @[Mux.scala 19:72:@32399.4]
  wire [7:0] _T_62679; // @[Mux.scala 19:72:@32406.4]
  wire [7:0] _T_62686; // @[Mux.scala 19:72:@32413.4]
  wire [15:0] _T_62687; // @[Mux.scala 19:72:@32414.4]
  wire [15:0] _T_62689; // @[Mux.scala 19:72:@32415.4]
  wire [7:0] _T_62696; // @[Mux.scala 19:72:@32422.4]
  wire [7:0] _T_62703; // @[Mux.scala 19:72:@32429.4]
  wire [15:0] _T_62704; // @[Mux.scala 19:72:@32430.4]
  wire [15:0] _T_62706; // @[Mux.scala 19:72:@32431.4]
  wire [7:0] _T_62713; // @[Mux.scala 19:72:@32438.4]
  wire [7:0] _T_62720; // @[Mux.scala 19:72:@32445.4]
  wire [15:0] _T_62721; // @[Mux.scala 19:72:@32446.4]
  wire [15:0] _T_62723; // @[Mux.scala 19:72:@32447.4]
  wire [7:0] _T_62730; // @[Mux.scala 19:72:@32454.4]
  wire [7:0] _T_62737; // @[Mux.scala 19:72:@32461.4]
  wire [15:0] _T_62738; // @[Mux.scala 19:72:@32462.4]
  wire [15:0] _T_62740; // @[Mux.scala 19:72:@32463.4]
  wire [7:0] _T_62747; // @[Mux.scala 19:72:@32470.4]
  wire [7:0] _T_62754; // @[Mux.scala 19:72:@32477.4]
  wire [15:0] _T_62755; // @[Mux.scala 19:72:@32478.4]
  wire [15:0] _T_62757; // @[Mux.scala 19:72:@32479.4]
  wire [15:0] _T_62772; // @[Mux.scala 19:72:@32494.4]
  wire [15:0] _T_62774; // @[Mux.scala 19:72:@32495.4]
  wire [15:0] _T_62789; // @[Mux.scala 19:72:@32510.4]
  wire [15:0] _T_62791; // @[Mux.scala 19:72:@32511.4]
  wire [15:0] _T_62806; // @[Mux.scala 19:72:@32526.4]
  wire [15:0] _T_62808; // @[Mux.scala 19:72:@32527.4]
  wire [15:0] _T_62823; // @[Mux.scala 19:72:@32542.4]
  wire [15:0] _T_62825; // @[Mux.scala 19:72:@32543.4]
  wire [15:0] _T_62840; // @[Mux.scala 19:72:@32558.4]
  wire [15:0] _T_62842; // @[Mux.scala 19:72:@32559.4]
  wire [15:0] _T_62857; // @[Mux.scala 19:72:@32574.4]
  wire [15:0] _T_62859; // @[Mux.scala 19:72:@32575.4]
  wire [15:0] _T_62874; // @[Mux.scala 19:72:@32590.4]
  wire [15:0] _T_62876; // @[Mux.scala 19:72:@32591.4]
  wire [15:0] _T_62891; // @[Mux.scala 19:72:@32606.4]
  wire [15:0] _T_62893; // @[Mux.scala 19:72:@32607.4]
  wire [15:0] _T_62894; // @[Mux.scala 19:72:@32608.4]
  wire [15:0] _T_62895; // @[Mux.scala 19:72:@32609.4]
  wire [15:0] _T_62896; // @[Mux.scala 19:72:@32610.4]
  wire [15:0] _T_62897; // @[Mux.scala 19:72:@32611.4]
  wire [15:0] _T_62898; // @[Mux.scala 19:72:@32612.4]
  wire [15:0] _T_62899; // @[Mux.scala 19:72:@32613.4]
  wire [15:0] _T_62900; // @[Mux.scala 19:72:@32614.4]
  wire [15:0] _T_62901; // @[Mux.scala 19:72:@32615.4]
  wire [15:0] _T_62902; // @[Mux.scala 19:72:@32616.4]
  wire [15:0] _T_62903; // @[Mux.scala 19:72:@32617.4]
  wire [15:0] _T_62904; // @[Mux.scala 19:72:@32618.4]
  wire [15:0] _T_62905; // @[Mux.scala 19:72:@32619.4]
  wire [15:0] _T_62906; // @[Mux.scala 19:72:@32620.4]
  wire [15:0] _T_62907; // @[Mux.scala 19:72:@32621.4]
  wire [15:0] _T_62908; // @[Mux.scala 19:72:@32622.4]
  wire [7:0] _T_63486; // @[Mux.scala 19:72:@32972.4]
  wire [7:0] _T_63493; // @[Mux.scala 19:72:@32979.4]
  wire [15:0] _T_63494; // @[Mux.scala 19:72:@32980.4]
  wire [15:0] _T_63496; // @[Mux.scala 19:72:@32981.4]
  wire [7:0] _T_63503; // @[Mux.scala 19:72:@32988.4]
  wire [7:0] _T_63510; // @[Mux.scala 19:72:@32995.4]
  wire [15:0] _T_63511; // @[Mux.scala 19:72:@32996.4]
  wire [15:0] _T_63513; // @[Mux.scala 19:72:@32997.4]
  wire [7:0] _T_63520; // @[Mux.scala 19:72:@33004.4]
  wire [7:0] _T_63527; // @[Mux.scala 19:72:@33011.4]
  wire [15:0] _T_63528; // @[Mux.scala 19:72:@33012.4]
  wire [15:0] _T_63530; // @[Mux.scala 19:72:@33013.4]
  wire [7:0] _T_63537; // @[Mux.scala 19:72:@33020.4]
  wire [7:0] _T_63544; // @[Mux.scala 19:72:@33027.4]
  wire [15:0] _T_63545; // @[Mux.scala 19:72:@33028.4]
  wire [15:0] _T_63547; // @[Mux.scala 19:72:@33029.4]
  wire [7:0] _T_63554; // @[Mux.scala 19:72:@33036.4]
  wire [7:0] _T_63561; // @[Mux.scala 19:72:@33043.4]
  wire [15:0] _T_63562; // @[Mux.scala 19:72:@33044.4]
  wire [15:0] _T_63564; // @[Mux.scala 19:72:@33045.4]
  wire [7:0] _T_63571; // @[Mux.scala 19:72:@33052.4]
  wire [7:0] _T_63578; // @[Mux.scala 19:72:@33059.4]
  wire [15:0] _T_63579; // @[Mux.scala 19:72:@33060.4]
  wire [15:0] _T_63581; // @[Mux.scala 19:72:@33061.4]
  wire [7:0] _T_63588; // @[Mux.scala 19:72:@33068.4]
  wire [7:0] _T_63595; // @[Mux.scala 19:72:@33075.4]
  wire [15:0] _T_63596; // @[Mux.scala 19:72:@33076.4]
  wire [15:0] _T_63598; // @[Mux.scala 19:72:@33077.4]
  wire [7:0] _T_63605; // @[Mux.scala 19:72:@33084.4]
  wire [7:0] _T_63612; // @[Mux.scala 19:72:@33091.4]
  wire [15:0] _T_63613; // @[Mux.scala 19:72:@33092.4]
  wire [15:0] _T_63615; // @[Mux.scala 19:72:@33093.4]
  wire [15:0] _T_63630; // @[Mux.scala 19:72:@33108.4]
  wire [15:0] _T_63632; // @[Mux.scala 19:72:@33109.4]
  wire [15:0] _T_63647; // @[Mux.scala 19:72:@33124.4]
  wire [15:0] _T_63649; // @[Mux.scala 19:72:@33125.4]
  wire [15:0] _T_63664; // @[Mux.scala 19:72:@33140.4]
  wire [15:0] _T_63666; // @[Mux.scala 19:72:@33141.4]
  wire [15:0] _T_63681; // @[Mux.scala 19:72:@33156.4]
  wire [15:0] _T_63683; // @[Mux.scala 19:72:@33157.4]
  wire [15:0] _T_63698; // @[Mux.scala 19:72:@33172.4]
  wire [15:0] _T_63700; // @[Mux.scala 19:72:@33173.4]
  wire [15:0] _T_63715; // @[Mux.scala 19:72:@33188.4]
  wire [15:0] _T_63717; // @[Mux.scala 19:72:@33189.4]
  wire [15:0] _T_63732; // @[Mux.scala 19:72:@33204.4]
  wire [15:0] _T_63734; // @[Mux.scala 19:72:@33205.4]
  wire [15:0] _T_63749; // @[Mux.scala 19:72:@33220.4]
  wire [15:0] _T_63751; // @[Mux.scala 19:72:@33221.4]
  wire [15:0] _T_63752; // @[Mux.scala 19:72:@33222.4]
  wire [15:0] _T_63753; // @[Mux.scala 19:72:@33223.4]
  wire [15:0] _T_63754; // @[Mux.scala 19:72:@33224.4]
  wire [15:0] _T_63755; // @[Mux.scala 19:72:@33225.4]
  wire [15:0] _T_63756; // @[Mux.scala 19:72:@33226.4]
  wire [15:0] _T_63757; // @[Mux.scala 19:72:@33227.4]
  wire [15:0] _T_63758; // @[Mux.scala 19:72:@33228.4]
  wire [15:0] _T_63759; // @[Mux.scala 19:72:@33229.4]
  wire [15:0] _T_63760; // @[Mux.scala 19:72:@33230.4]
  wire [15:0] _T_63761; // @[Mux.scala 19:72:@33231.4]
  wire [15:0] _T_63762; // @[Mux.scala 19:72:@33232.4]
  wire [15:0] _T_63763; // @[Mux.scala 19:72:@33233.4]
  wire [15:0] _T_63764; // @[Mux.scala 19:72:@33234.4]
  wire [15:0] _T_63765; // @[Mux.scala 19:72:@33235.4]
  wire [15:0] _T_63766; // @[Mux.scala 19:72:@33236.4]
  wire [7:0] _T_64344; // @[Mux.scala 19:72:@33586.4]
  wire [7:0] _T_64351; // @[Mux.scala 19:72:@33593.4]
  wire [15:0] _T_64352; // @[Mux.scala 19:72:@33594.4]
  wire [15:0] _T_64354; // @[Mux.scala 19:72:@33595.4]
  wire [7:0] _T_64361; // @[Mux.scala 19:72:@33602.4]
  wire [7:0] _T_64368; // @[Mux.scala 19:72:@33609.4]
  wire [15:0] _T_64369; // @[Mux.scala 19:72:@33610.4]
  wire [15:0] _T_64371; // @[Mux.scala 19:72:@33611.4]
  wire [7:0] _T_64378; // @[Mux.scala 19:72:@33618.4]
  wire [7:0] _T_64385; // @[Mux.scala 19:72:@33625.4]
  wire [15:0] _T_64386; // @[Mux.scala 19:72:@33626.4]
  wire [15:0] _T_64388; // @[Mux.scala 19:72:@33627.4]
  wire [7:0] _T_64395; // @[Mux.scala 19:72:@33634.4]
  wire [7:0] _T_64402; // @[Mux.scala 19:72:@33641.4]
  wire [15:0] _T_64403; // @[Mux.scala 19:72:@33642.4]
  wire [15:0] _T_64405; // @[Mux.scala 19:72:@33643.4]
  wire [7:0] _T_64412; // @[Mux.scala 19:72:@33650.4]
  wire [7:0] _T_64419; // @[Mux.scala 19:72:@33657.4]
  wire [15:0] _T_64420; // @[Mux.scala 19:72:@33658.4]
  wire [15:0] _T_64422; // @[Mux.scala 19:72:@33659.4]
  wire [7:0] _T_64429; // @[Mux.scala 19:72:@33666.4]
  wire [7:0] _T_64436; // @[Mux.scala 19:72:@33673.4]
  wire [15:0] _T_64437; // @[Mux.scala 19:72:@33674.4]
  wire [15:0] _T_64439; // @[Mux.scala 19:72:@33675.4]
  wire [7:0] _T_64446; // @[Mux.scala 19:72:@33682.4]
  wire [7:0] _T_64453; // @[Mux.scala 19:72:@33689.4]
  wire [15:0] _T_64454; // @[Mux.scala 19:72:@33690.4]
  wire [15:0] _T_64456; // @[Mux.scala 19:72:@33691.4]
  wire [7:0] _T_64463; // @[Mux.scala 19:72:@33698.4]
  wire [7:0] _T_64470; // @[Mux.scala 19:72:@33705.4]
  wire [15:0] _T_64471; // @[Mux.scala 19:72:@33706.4]
  wire [15:0] _T_64473; // @[Mux.scala 19:72:@33707.4]
  wire [15:0] _T_64488; // @[Mux.scala 19:72:@33722.4]
  wire [15:0] _T_64490; // @[Mux.scala 19:72:@33723.4]
  wire [15:0] _T_64505; // @[Mux.scala 19:72:@33738.4]
  wire [15:0] _T_64507; // @[Mux.scala 19:72:@33739.4]
  wire [15:0] _T_64522; // @[Mux.scala 19:72:@33754.4]
  wire [15:0] _T_64524; // @[Mux.scala 19:72:@33755.4]
  wire [15:0] _T_64539; // @[Mux.scala 19:72:@33770.4]
  wire [15:0] _T_64541; // @[Mux.scala 19:72:@33771.4]
  wire [15:0] _T_64556; // @[Mux.scala 19:72:@33786.4]
  wire [15:0] _T_64558; // @[Mux.scala 19:72:@33787.4]
  wire [15:0] _T_64573; // @[Mux.scala 19:72:@33802.4]
  wire [15:0] _T_64575; // @[Mux.scala 19:72:@33803.4]
  wire [15:0] _T_64590; // @[Mux.scala 19:72:@33818.4]
  wire [15:0] _T_64592; // @[Mux.scala 19:72:@33819.4]
  wire [15:0] _T_64607; // @[Mux.scala 19:72:@33834.4]
  wire [15:0] _T_64609; // @[Mux.scala 19:72:@33835.4]
  wire [15:0] _T_64610; // @[Mux.scala 19:72:@33836.4]
  wire [15:0] _T_64611; // @[Mux.scala 19:72:@33837.4]
  wire [15:0] _T_64612; // @[Mux.scala 19:72:@33838.4]
  wire [15:0] _T_64613; // @[Mux.scala 19:72:@33839.4]
  wire [15:0] _T_64614; // @[Mux.scala 19:72:@33840.4]
  wire [15:0] _T_64615; // @[Mux.scala 19:72:@33841.4]
  wire [15:0] _T_64616; // @[Mux.scala 19:72:@33842.4]
  wire [15:0] _T_64617; // @[Mux.scala 19:72:@33843.4]
  wire [15:0] _T_64618; // @[Mux.scala 19:72:@33844.4]
  wire [15:0] _T_64619; // @[Mux.scala 19:72:@33845.4]
  wire [15:0] _T_64620; // @[Mux.scala 19:72:@33846.4]
  wire [15:0] _T_64621; // @[Mux.scala 19:72:@33847.4]
  wire [15:0] _T_64622; // @[Mux.scala 19:72:@33848.4]
  wire [15:0] _T_64623; // @[Mux.scala 19:72:@33849.4]
  wire [15:0] _T_64624; // @[Mux.scala 19:72:@33850.4]
  wire [7:0] _T_65202; // @[Mux.scala 19:72:@34200.4]
  wire [7:0] _T_65209; // @[Mux.scala 19:72:@34207.4]
  wire [15:0] _T_65210; // @[Mux.scala 19:72:@34208.4]
  wire [15:0] _T_65212; // @[Mux.scala 19:72:@34209.4]
  wire [7:0] _T_65219; // @[Mux.scala 19:72:@34216.4]
  wire [7:0] _T_65226; // @[Mux.scala 19:72:@34223.4]
  wire [15:0] _T_65227; // @[Mux.scala 19:72:@34224.4]
  wire [15:0] _T_65229; // @[Mux.scala 19:72:@34225.4]
  wire [7:0] _T_65236; // @[Mux.scala 19:72:@34232.4]
  wire [7:0] _T_65243; // @[Mux.scala 19:72:@34239.4]
  wire [15:0] _T_65244; // @[Mux.scala 19:72:@34240.4]
  wire [15:0] _T_65246; // @[Mux.scala 19:72:@34241.4]
  wire [7:0] _T_65253; // @[Mux.scala 19:72:@34248.4]
  wire [7:0] _T_65260; // @[Mux.scala 19:72:@34255.4]
  wire [15:0] _T_65261; // @[Mux.scala 19:72:@34256.4]
  wire [15:0] _T_65263; // @[Mux.scala 19:72:@34257.4]
  wire [7:0] _T_65270; // @[Mux.scala 19:72:@34264.4]
  wire [7:0] _T_65277; // @[Mux.scala 19:72:@34271.4]
  wire [15:0] _T_65278; // @[Mux.scala 19:72:@34272.4]
  wire [15:0] _T_65280; // @[Mux.scala 19:72:@34273.4]
  wire [7:0] _T_65287; // @[Mux.scala 19:72:@34280.4]
  wire [7:0] _T_65294; // @[Mux.scala 19:72:@34287.4]
  wire [15:0] _T_65295; // @[Mux.scala 19:72:@34288.4]
  wire [15:0] _T_65297; // @[Mux.scala 19:72:@34289.4]
  wire [7:0] _T_65304; // @[Mux.scala 19:72:@34296.4]
  wire [7:0] _T_65311; // @[Mux.scala 19:72:@34303.4]
  wire [15:0] _T_65312; // @[Mux.scala 19:72:@34304.4]
  wire [15:0] _T_65314; // @[Mux.scala 19:72:@34305.4]
  wire [7:0] _T_65321; // @[Mux.scala 19:72:@34312.4]
  wire [7:0] _T_65328; // @[Mux.scala 19:72:@34319.4]
  wire [15:0] _T_65329; // @[Mux.scala 19:72:@34320.4]
  wire [15:0] _T_65331; // @[Mux.scala 19:72:@34321.4]
  wire [15:0] _T_65346; // @[Mux.scala 19:72:@34336.4]
  wire [15:0] _T_65348; // @[Mux.scala 19:72:@34337.4]
  wire [15:0] _T_65363; // @[Mux.scala 19:72:@34352.4]
  wire [15:0] _T_65365; // @[Mux.scala 19:72:@34353.4]
  wire [15:0] _T_65380; // @[Mux.scala 19:72:@34368.4]
  wire [15:0] _T_65382; // @[Mux.scala 19:72:@34369.4]
  wire [15:0] _T_65397; // @[Mux.scala 19:72:@34384.4]
  wire [15:0] _T_65399; // @[Mux.scala 19:72:@34385.4]
  wire [15:0] _T_65414; // @[Mux.scala 19:72:@34400.4]
  wire [15:0] _T_65416; // @[Mux.scala 19:72:@34401.4]
  wire [15:0] _T_65431; // @[Mux.scala 19:72:@34416.4]
  wire [15:0] _T_65433; // @[Mux.scala 19:72:@34417.4]
  wire [15:0] _T_65448; // @[Mux.scala 19:72:@34432.4]
  wire [15:0] _T_65450; // @[Mux.scala 19:72:@34433.4]
  wire [15:0] _T_65465; // @[Mux.scala 19:72:@34448.4]
  wire [15:0] _T_65467; // @[Mux.scala 19:72:@34449.4]
  wire [15:0] _T_65468; // @[Mux.scala 19:72:@34450.4]
  wire [15:0] _T_65469; // @[Mux.scala 19:72:@34451.4]
  wire [15:0] _T_65470; // @[Mux.scala 19:72:@34452.4]
  wire [15:0] _T_65471; // @[Mux.scala 19:72:@34453.4]
  wire [15:0] _T_65472; // @[Mux.scala 19:72:@34454.4]
  wire [15:0] _T_65473; // @[Mux.scala 19:72:@34455.4]
  wire [15:0] _T_65474; // @[Mux.scala 19:72:@34456.4]
  wire [15:0] _T_65475; // @[Mux.scala 19:72:@34457.4]
  wire [15:0] _T_65476; // @[Mux.scala 19:72:@34458.4]
  wire [15:0] _T_65477; // @[Mux.scala 19:72:@34459.4]
  wire [15:0] _T_65478; // @[Mux.scala 19:72:@34460.4]
  wire [15:0] _T_65479; // @[Mux.scala 19:72:@34461.4]
  wire [15:0] _T_65480; // @[Mux.scala 19:72:@34462.4]
  wire [15:0] _T_65481; // @[Mux.scala 19:72:@34463.4]
  wire [15:0] _T_65482; // @[Mux.scala 19:72:@34464.4]
  reg  storeAddrNotKnownFlagsPReg_0_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_419;
  reg  storeAddrNotKnownFlagsPReg_0_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_420;
  reg  storeAddrNotKnownFlagsPReg_0_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_421;
  reg  storeAddrNotKnownFlagsPReg_0_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_422;
  reg  storeAddrNotKnownFlagsPReg_0_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_423;
  reg  storeAddrNotKnownFlagsPReg_0_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_424;
  reg  storeAddrNotKnownFlagsPReg_0_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_425;
  reg  storeAddrNotKnownFlagsPReg_0_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_426;
  reg  storeAddrNotKnownFlagsPReg_0_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_427;
  reg  storeAddrNotKnownFlagsPReg_0_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_428;
  reg  storeAddrNotKnownFlagsPReg_0_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_429;
  reg  storeAddrNotKnownFlagsPReg_0_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_430;
  reg  storeAddrNotKnownFlagsPReg_0_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_431;
  reg  storeAddrNotKnownFlagsPReg_0_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_432;
  reg  storeAddrNotKnownFlagsPReg_0_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_433;
  reg  storeAddrNotKnownFlagsPReg_0_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_434;
  reg  storeAddrNotKnownFlagsPReg_1_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_435;
  reg  storeAddrNotKnownFlagsPReg_1_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_436;
  reg  storeAddrNotKnownFlagsPReg_1_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_437;
  reg  storeAddrNotKnownFlagsPReg_1_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_438;
  reg  storeAddrNotKnownFlagsPReg_1_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_439;
  reg  storeAddrNotKnownFlagsPReg_1_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_440;
  reg  storeAddrNotKnownFlagsPReg_1_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_441;
  reg  storeAddrNotKnownFlagsPReg_1_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_442;
  reg  storeAddrNotKnownFlagsPReg_1_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_443;
  reg  storeAddrNotKnownFlagsPReg_1_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_444;
  reg  storeAddrNotKnownFlagsPReg_1_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_445;
  reg  storeAddrNotKnownFlagsPReg_1_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_446;
  reg  storeAddrNotKnownFlagsPReg_1_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_447;
  reg  storeAddrNotKnownFlagsPReg_1_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_448;
  reg  storeAddrNotKnownFlagsPReg_1_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_449;
  reg  storeAddrNotKnownFlagsPReg_1_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_450;
  reg  storeAddrNotKnownFlagsPReg_2_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_451;
  reg  storeAddrNotKnownFlagsPReg_2_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_452;
  reg  storeAddrNotKnownFlagsPReg_2_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_453;
  reg  storeAddrNotKnownFlagsPReg_2_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_454;
  reg  storeAddrNotKnownFlagsPReg_2_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_455;
  reg  storeAddrNotKnownFlagsPReg_2_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_456;
  reg  storeAddrNotKnownFlagsPReg_2_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_457;
  reg  storeAddrNotKnownFlagsPReg_2_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_458;
  reg  storeAddrNotKnownFlagsPReg_2_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_459;
  reg  storeAddrNotKnownFlagsPReg_2_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_460;
  reg  storeAddrNotKnownFlagsPReg_2_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_461;
  reg  storeAddrNotKnownFlagsPReg_2_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_462;
  reg  storeAddrNotKnownFlagsPReg_2_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_463;
  reg  storeAddrNotKnownFlagsPReg_2_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_464;
  reg  storeAddrNotKnownFlagsPReg_2_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_465;
  reg  storeAddrNotKnownFlagsPReg_2_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_466;
  reg  storeAddrNotKnownFlagsPReg_3_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_467;
  reg  storeAddrNotKnownFlagsPReg_3_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_468;
  reg  storeAddrNotKnownFlagsPReg_3_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_469;
  reg  storeAddrNotKnownFlagsPReg_3_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_470;
  reg  storeAddrNotKnownFlagsPReg_3_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_471;
  reg  storeAddrNotKnownFlagsPReg_3_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_472;
  reg  storeAddrNotKnownFlagsPReg_3_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_473;
  reg  storeAddrNotKnownFlagsPReg_3_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_474;
  reg  storeAddrNotKnownFlagsPReg_3_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_475;
  reg  storeAddrNotKnownFlagsPReg_3_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_476;
  reg  storeAddrNotKnownFlagsPReg_3_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_477;
  reg  storeAddrNotKnownFlagsPReg_3_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_478;
  reg  storeAddrNotKnownFlagsPReg_3_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_479;
  reg  storeAddrNotKnownFlagsPReg_3_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_480;
  reg  storeAddrNotKnownFlagsPReg_3_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_481;
  reg  storeAddrNotKnownFlagsPReg_3_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_482;
  reg  storeAddrNotKnownFlagsPReg_4_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_483;
  reg  storeAddrNotKnownFlagsPReg_4_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_484;
  reg  storeAddrNotKnownFlagsPReg_4_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_485;
  reg  storeAddrNotKnownFlagsPReg_4_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_486;
  reg  storeAddrNotKnownFlagsPReg_4_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_487;
  reg  storeAddrNotKnownFlagsPReg_4_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_488;
  reg  storeAddrNotKnownFlagsPReg_4_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_489;
  reg  storeAddrNotKnownFlagsPReg_4_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_490;
  reg  storeAddrNotKnownFlagsPReg_4_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_491;
  reg  storeAddrNotKnownFlagsPReg_4_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_492;
  reg  storeAddrNotKnownFlagsPReg_4_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_493;
  reg  storeAddrNotKnownFlagsPReg_4_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_494;
  reg  storeAddrNotKnownFlagsPReg_4_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_495;
  reg  storeAddrNotKnownFlagsPReg_4_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_496;
  reg  storeAddrNotKnownFlagsPReg_4_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_497;
  reg  storeAddrNotKnownFlagsPReg_4_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_498;
  reg  storeAddrNotKnownFlagsPReg_5_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_499;
  reg  storeAddrNotKnownFlagsPReg_5_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_500;
  reg  storeAddrNotKnownFlagsPReg_5_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_501;
  reg  storeAddrNotKnownFlagsPReg_5_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_502;
  reg  storeAddrNotKnownFlagsPReg_5_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_503;
  reg  storeAddrNotKnownFlagsPReg_5_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_504;
  reg  storeAddrNotKnownFlagsPReg_5_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_505;
  reg  storeAddrNotKnownFlagsPReg_5_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_506;
  reg  storeAddrNotKnownFlagsPReg_5_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_507;
  reg  storeAddrNotKnownFlagsPReg_5_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_508;
  reg  storeAddrNotKnownFlagsPReg_5_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_509;
  reg  storeAddrNotKnownFlagsPReg_5_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_510;
  reg  storeAddrNotKnownFlagsPReg_5_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_511;
  reg  storeAddrNotKnownFlagsPReg_5_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_512;
  reg  storeAddrNotKnownFlagsPReg_5_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_513;
  reg  storeAddrNotKnownFlagsPReg_5_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_514;
  reg  storeAddrNotKnownFlagsPReg_6_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_515;
  reg  storeAddrNotKnownFlagsPReg_6_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_516;
  reg  storeAddrNotKnownFlagsPReg_6_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_517;
  reg  storeAddrNotKnownFlagsPReg_6_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_518;
  reg  storeAddrNotKnownFlagsPReg_6_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_519;
  reg  storeAddrNotKnownFlagsPReg_6_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_520;
  reg  storeAddrNotKnownFlagsPReg_6_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_521;
  reg  storeAddrNotKnownFlagsPReg_6_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_522;
  reg  storeAddrNotKnownFlagsPReg_6_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_523;
  reg  storeAddrNotKnownFlagsPReg_6_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_524;
  reg  storeAddrNotKnownFlagsPReg_6_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_525;
  reg  storeAddrNotKnownFlagsPReg_6_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_526;
  reg  storeAddrNotKnownFlagsPReg_6_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_527;
  reg  storeAddrNotKnownFlagsPReg_6_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_528;
  reg  storeAddrNotKnownFlagsPReg_6_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_529;
  reg  storeAddrNotKnownFlagsPReg_6_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_530;
  reg  storeAddrNotKnownFlagsPReg_7_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_531;
  reg  storeAddrNotKnownFlagsPReg_7_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_532;
  reg  storeAddrNotKnownFlagsPReg_7_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_533;
  reg  storeAddrNotKnownFlagsPReg_7_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_534;
  reg  storeAddrNotKnownFlagsPReg_7_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_535;
  reg  storeAddrNotKnownFlagsPReg_7_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_536;
  reg  storeAddrNotKnownFlagsPReg_7_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_537;
  reg  storeAddrNotKnownFlagsPReg_7_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_538;
  reg  storeAddrNotKnownFlagsPReg_7_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_539;
  reg  storeAddrNotKnownFlagsPReg_7_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_540;
  reg  storeAddrNotKnownFlagsPReg_7_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_541;
  reg  storeAddrNotKnownFlagsPReg_7_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_542;
  reg  storeAddrNotKnownFlagsPReg_7_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_543;
  reg  storeAddrNotKnownFlagsPReg_7_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_544;
  reg  storeAddrNotKnownFlagsPReg_7_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_545;
  reg  storeAddrNotKnownFlagsPReg_7_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_546;
  reg  storeAddrNotKnownFlagsPReg_8_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_547;
  reg  storeAddrNotKnownFlagsPReg_8_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_548;
  reg  storeAddrNotKnownFlagsPReg_8_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_549;
  reg  storeAddrNotKnownFlagsPReg_8_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_550;
  reg  storeAddrNotKnownFlagsPReg_8_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_551;
  reg  storeAddrNotKnownFlagsPReg_8_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_552;
  reg  storeAddrNotKnownFlagsPReg_8_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_553;
  reg  storeAddrNotKnownFlagsPReg_8_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_554;
  reg  storeAddrNotKnownFlagsPReg_8_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_555;
  reg  storeAddrNotKnownFlagsPReg_8_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_556;
  reg  storeAddrNotKnownFlagsPReg_8_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_557;
  reg  storeAddrNotKnownFlagsPReg_8_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_558;
  reg  storeAddrNotKnownFlagsPReg_8_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_559;
  reg  storeAddrNotKnownFlagsPReg_8_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_560;
  reg  storeAddrNotKnownFlagsPReg_8_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_561;
  reg  storeAddrNotKnownFlagsPReg_8_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_562;
  reg  storeAddrNotKnownFlagsPReg_9_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_563;
  reg  storeAddrNotKnownFlagsPReg_9_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_564;
  reg  storeAddrNotKnownFlagsPReg_9_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_565;
  reg  storeAddrNotKnownFlagsPReg_9_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_566;
  reg  storeAddrNotKnownFlagsPReg_9_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_567;
  reg  storeAddrNotKnownFlagsPReg_9_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_568;
  reg  storeAddrNotKnownFlagsPReg_9_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_569;
  reg  storeAddrNotKnownFlagsPReg_9_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_570;
  reg  storeAddrNotKnownFlagsPReg_9_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_571;
  reg  storeAddrNotKnownFlagsPReg_9_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_572;
  reg  storeAddrNotKnownFlagsPReg_9_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_573;
  reg  storeAddrNotKnownFlagsPReg_9_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_574;
  reg  storeAddrNotKnownFlagsPReg_9_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_575;
  reg  storeAddrNotKnownFlagsPReg_9_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_576;
  reg  storeAddrNotKnownFlagsPReg_9_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_577;
  reg  storeAddrNotKnownFlagsPReg_9_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_578;
  reg  storeAddrNotKnownFlagsPReg_10_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_579;
  reg  storeAddrNotKnownFlagsPReg_10_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_580;
  reg  storeAddrNotKnownFlagsPReg_10_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_581;
  reg  storeAddrNotKnownFlagsPReg_10_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_582;
  reg  storeAddrNotKnownFlagsPReg_10_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_583;
  reg  storeAddrNotKnownFlagsPReg_10_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_584;
  reg  storeAddrNotKnownFlagsPReg_10_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_585;
  reg  storeAddrNotKnownFlagsPReg_10_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_586;
  reg  storeAddrNotKnownFlagsPReg_10_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_587;
  reg  storeAddrNotKnownFlagsPReg_10_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_588;
  reg  storeAddrNotKnownFlagsPReg_10_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_589;
  reg  storeAddrNotKnownFlagsPReg_10_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_590;
  reg  storeAddrNotKnownFlagsPReg_10_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_591;
  reg  storeAddrNotKnownFlagsPReg_10_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_592;
  reg  storeAddrNotKnownFlagsPReg_10_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_593;
  reg  storeAddrNotKnownFlagsPReg_10_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_594;
  reg  storeAddrNotKnownFlagsPReg_11_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_595;
  reg  storeAddrNotKnownFlagsPReg_11_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_596;
  reg  storeAddrNotKnownFlagsPReg_11_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_597;
  reg  storeAddrNotKnownFlagsPReg_11_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_598;
  reg  storeAddrNotKnownFlagsPReg_11_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_599;
  reg  storeAddrNotKnownFlagsPReg_11_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_600;
  reg  storeAddrNotKnownFlagsPReg_11_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_601;
  reg  storeAddrNotKnownFlagsPReg_11_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_602;
  reg  storeAddrNotKnownFlagsPReg_11_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_603;
  reg  storeAddrNotKnownFlagsPReg_11_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_604;
  reg  storeAddrNotKnownFlagsPReg_11_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_605;
  reg  storeAddrNotKnownFlagsPReg_11_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_606;
  reg  storeAddrNotKnownFlagsPReg_11_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_607;
  reg  storeAddrNotKnownFlagsPReg_11_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_608;
  reg  storeAddrNotKnownFlagsPReg_11_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_609;
  reg  storeAddrNotKnownFlagsPReg_11_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_610;
  reg  storeAddrNotKnownFlagsPReg_12_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_611;
  reg  storeAddrNotKnownFlagsPReg_12_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_612;
  reg  storeAddrNotKnownFlagsPReg_12_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_613;
  reg  storeAddrNotKnownFlagsPReg_12_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_614;
  reg  storeAddrNotKnownFlagsPReg_12_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_615;
  reg  storeAddrNotKnownFlagsPReg_12_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_616;
  reg  storeAddrNotKnownFlagsPReg_12_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_617;
  reg  storeAddrNotKnownFlagsPReg_12_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_618;
  reg  storeAddrNotKnownFlagsPReg_12_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_619;
  reg  storeAddrNotKnownFlagsPReg_12_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_620;
  reg  storeAddrNotKnownFlagsPReg_12_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_621;
  reg  storeAddrNotKnownFlagsPReg_12_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_622;
  reg  storeAddrNotKnownFlagsPReg_12_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_623;
  reg  storeAddrNotKnownFlagsPReg_12_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_624;
  reg  storeAddrNotKnownFlagsPReg_12_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_625;
  reg  storeAddrNotKnownFlagsPReg_12_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_626;
  reg  storeAddrNotKnownFlagsPReg_13_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_627;
  reg  storeAddrNotKnownFlagsPReg_13_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_628;
  reg  storeAddrNotKnownFlagsPReg_13_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_629;
  reg  storeAddrNotKnownFlagsPReg_13_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_630;
  reg  storeAddrNotKnownFlagsPReg_13_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_631;
  reg  storeAddrNotKnownFlagsPReg_13_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_632;
  reg  storeAddrNotKnownFlagsPReg_13_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_633;
  reg  storeAddrNotKnownFlagsPReg_13_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_634;
  reg  storeAddrNotKnownFlagsPReg_13_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_635;
  reg  storeAddrNotKnownFlagsPReg_13_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_636;
  reg  storeAddrNotKnownFlagsPReg_13_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_637;
  reg  storeAddrNotKnownFlagsPReg_13_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_638;
  reg  storeAddrNotKnownFlagsPReg_13_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_639;
  reg  storeAddrNotKnownFlagsPReg_13_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_640;
  reg  storeAddrNotKnownFlagsPReg_13_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_641;
  reg  storeAddrNotKnownFlagsPReg_13_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_642;
  reg  storeAddrNotKnownFlagsPReg_14_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_643;
  reg  storeAddrNotKnownFlagsPReg_14_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_644;
  reg  storeAddrNotKnownFlagsPReg_14_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_645;
  reg  storeAddrNotKnownFlagsPReg_14_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_646;
  reg  storeAddrNotKnownFlagsPReg_14_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_647;
  reg  storeAddrNotKnownFlagsPReg_14_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_648;
  reg  storeAddrNotKnownFlagsPReg_14_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_649;
  reg  storeAddrNotKnownFlagsPReg_14_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_650;
  reg  storeAddrNotKnownFlagsPReg_14_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_651;
  reg  storeAddrNotKnownFlagsPReg_14_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_652;
  reg  storeAddrNotKnownFlagsPReg_14_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_653;
  reg  storeAddrNotKnownFlagsPReg_14_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_654;
  reg  storeAddrNotKnownFlagsPReg_14_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_655;
  reg  storeAddrNotKnownFlagsPReg_14_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_656;
  reg  storeAddrNotKnownFlagsPReg_14_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_657;
  reg  storeAddrNotKnownFlagsPReg_14_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_658;
  reg  storeAddrNotKnownFlagsPReg_15_0; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_659;
  reg  storeAddrNotKnownFlagsPReg_15_1; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_660;
  reg  storeAddrNotKnownFlagsPReg_15_2; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_661;
  reg  storeAddrNotKnownFlagsPReg_15_3; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_662;
  reg  storeAddrNotKnownFlagsPReg_15_4; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_663;
  reg  storeAddrNotKnownFlagsPReg_15_5; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_664;
  reg  storeAddrNotKnownFlagsPReg_15_6; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_665;
  reg  storeAddrNotKnownFlagsPReg_15_7; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_666;
  reg  storeAddrNotKnownFlagsPReg_15_8; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_667;
  reg  storeAddrNotKnownFlagsPReg_15_9; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_668;
  reg  storeAddrNotKnownFlagsPReg_15_10; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_669;
  reg  storeAddrNotKnownFlagsPReg_15_11; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_670;
  reg  storeAddrNotKnownFlagsPReg_15_12; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_671;
  reg  storeAddrNotKnownFlagsPReg_15_13; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_672;
  reg  storeAddrNotKnownFlagsPReg_15_14; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_673;
  reg  storeAddrNotKnownFlagsPReg_15_15; // @[AxiLoadQueue.scala 167:43:@34757.4]
  reg [31:0] _RAND_674;
  reg  shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_675;
  reg  shiftedStoreDataKnownPReg_1; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_676;
  reg  shiftedStoreDataKnownPReg_2; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_677;
  reg  shiftedStoreDataKnownPReg_3; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_678;
  reg  shiftedStoreDataKnownPReg_4; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_679;
  reg  shiftedStoreDataKnownPReg_5; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_680;
  reg  shiftedStoreDataKnownPReg_6; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_681;
  reg  shiftedStoreDataKnownPReg_7; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_682;
  reg  shiftedStoreDataKnownPReg_8; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_683;
  reg  shiftedStoreDataKnownPReg_9; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_684;
  reg  shiftedStoreDataKnownPReg_10; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_685;
  reg  shiftedStoreDataKnownPReg_11; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_686;
  reg  shiftedStoreDataKnownPReg_12; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_687;
  reg  shiftedStoreDataKnownPReg_13; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_688;
  reg  shiftedStoreDataKnownPReg_14; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_689;
  reg  shiftedStoreDataKnownPReg_15; // @[AxiLoadQueue.scala 168:42:@35014.4]
  reg [31:0] _RAND_690;
  reg [31:0] shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_691;
  reg [31:0] shiftedStoreDataQPreg_1; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_692;
  reg [31:0] shiftedStoreDataQPreg_2; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_693;
  reg [31:0] shiftedStoreDataQPreg_3; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_694;
  reg [31:0] shiftedStoreDataQPreg_4; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_695;
  reg [31:0] shiftedStoreDataQPreg_5; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_696;
  reg [31:0] shiftedStoreDataQPreg_6; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_697;
  reg [31:0] shiftedStoreDataQPreg_7; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_698;
  reg [31:0] shiftedStoreDataQPreg_8; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_699;
  reg [31:0] shiftedStoreDataQPreg_9; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_700;
  reg [31:0] shiftedStoreDataQPreg_10; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_701;
  reg [31:0] shiftedStoreDataQPreg_11; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_702;
  reg [31:0] shiftedStoreDataQPreg_12; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_703;
  reg [31:0] shiftedStoreDataQPreg_13; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_704;
  reg [31:0] shiftedStoreDataQPreg_14; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_705;
  reg [31:0] shiftedStoreDataQPreg_15; // @[AxiLoadQueue.scala 169:38:@35031.4]
  reg [31:0] _RAND_706;
  reg  addrKnownPReg_0; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_707;
  reg  addrKnownPReg_1; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_708;
  reg  addrKnownPReg_2; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_709;
  reg  addrKnownPReg_3; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_710;
  reg  addrKnownPReg_4; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_711;
  reg  addrKnownPReg_5; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_712;
  reg  addrKnownPReg_6; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_713;
  reg  addrKnownPReg_7; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_714;
  reg  addrKnownPReg_8; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_715;
  reg  addrKnownPReg_9; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_716;
  reg  addrKnownPReg_10; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_717;
  reg  addrKnownPReg_11; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_718;
  reg  addrKnownPReg_12; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_719;
  reg  addrKnownPReg_13; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_720;
  reg  addrKnownPReg_14; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_721;
  reg  addrKnownPReg_15; // @[AxiLoadQueue.scala 170:30:@35048.4]
  reg [31:0] _RAND_722;
  reg  dataKnownPReg_0; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_723;
  reg  dataKnownPReg_1; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_724;
  reg  dataKnownPReg_2; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_725;
  reg  dataKnownPReg_3; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_726;
  reg  dataKnownPReg_4; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_727;
  reg  dataKnownPReg_5; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_728;
  reg  dataKnownPReg_6; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_729;
  reg  dataKnownPReg_7; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_730;
  reg  dataKnownPReg_8; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_731;
  reg  dataKnownPReg_9; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_732;
  reg  dataKnownPReg_10; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_733;
  reg  dataKnownPReg_11; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_734;
  reg  dataKnownPReg_12; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_735;
  reg  dataKnownPReg_13; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_736;
  reg  dataKnownPReg_14; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_737;
  reg  dataKnownPReg_15; // @[AxiLoadQueue.scala 171:30:@35065.4]
  reg [31:0] _RAND_738;
  wire [1:0] _T_88274; // @[AxiLoadQueue.scala 191:60:@35137.4]
  wire [1:0] _T_88275; // @[AxiLoadQueue.scala 191:60:@35138.4]
  wire [2:0] _T_88276; // @[AxiLoadQueue.scala 191:60:@35139.4]
  wire [2:0] _T_88277; // @[AxiLoadQueue.scala 191:60:@35140.4]
  wire [2:0] _T_88278; // @[AxiLoadQueue.scala 191:60:@35141.4]
  wire [2:0] _T_88279; // @[AxiLoadQueue.scala 191:60:@35142.4]
  wire [3:0] _T_88280; // @[AxiLoadQueue.scala 191:60:@35143.4]
  wire [3:0] _T_88281; // @[AxiLoadQueue.scala 191:60:@35144.4]
  wire [3:0] _T_88282; // @[AxiLoadQueue.scala 191:60:@35145.4]
  wire [3:0] _T_88283; // @[AxiLoadQueue.scala 191:60:@35146.4]
  wire [3:0] _T_88284; // @[AxiLoadQueue.scala 191:60:@35147.4]
  wire [3:0] _T_88285; // @[AxiLoadQueue.scala 191:60:@35148.4]
  wire [3:0] _T_88286; // @[AxiLoadQueue.scala 191:60:@35149.4]
  wire [3:0] _T_88287; // @[AxiLoadQueue.scala 191:60:@35150.4]
  wire  _T_88290; // @[AxiLoadQueue.scala 192:43:@35152.4]
  wire  _T_88291; // @[AxiLoadQueue.scala 192:43:@35153.4]
  wire  _T_88292; // @[AxiLoadQueue.scala 192:43:@35154.4]
  wire  _T_88293; // @[AxiLoadQueue.scala 192:43:@35155.4]
  wire  _T_88294; // @[AxiLoadQueue.scala 192:43:@35156.4]
  wire  _T_88295; // @[AxiLoadQueue.scala 192:43:@35157.4]
  wire  _T_88296; // @[AxiLoadQueue.scala 192:43:@35158.4]
  wire  _T_88297; // @[AxiLoadQueue.scala 192:43:@35159.4]
  wire  _T_88298; // @[AxiLoadQueue.scala 192:43:@35160.4]
  wire  _T_88299; // @[AxiLoadQueue.scala 192:43:@35161.4]
  wire  _T_88300; // @[AxiLoadQueue.scala 192:43:@35162.4]
  wire  _T_88301; // @[AxiLoadQueue.scala 192:43:@35163.4]
  wire  _T_88302; // @[AxiLoadQueue.scala 192:43:@35164.4]
  wire  _T_88303; // @[AxiLoadQueue.scala 192:43:@35165.4]
  wire  _T_88304; // @[AxiLoadQueue.scala 192:43:@35166.4]
  wire  _GEN_864; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_865; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_866; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_867; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_868; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_869; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_870; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_871; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_872; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_873; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_874; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_875; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_876; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_877; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_878; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_879; // @[AxiLoadQueue.scala 193:43:@35168.6]
  wire  _GEN_881; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_882; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_883; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_884; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_885; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_886; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_887; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_888; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_889; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_890; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_891; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_892; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_893; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_894; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire  _GEN_895; // @[AxiLoadQueue.scala 194:31:@35169.6]
  wire [31:0] _GEN_897; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_898; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_899; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_900; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_901; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_902; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_903; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_904; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_905; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_906; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_907; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_908; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_909; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_910; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire [31:0] _GEN_911; // @[AxiLoadQueue.scala 195:31:@35170.6]
  wire  lastConflict_0_0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_1; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_2; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_3; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_4; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_5; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_6; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_7; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_8; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_9; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_10; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_11; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_12; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_13; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_14; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  lastConflict_0_15; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire  canBypass_0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire [31:0] bypassVal_0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  wire [1:0] _T_88410; // @[AxiLoadQueue.scala 191:60:@35224.4]
  wire [1:0] _T_88411; // @[AxiLoadQueue.scala 191:60:@35225.4]
  wire [2:0] _T_88412; // @[AxiLoadQueue.scala 191:60:@35226.4]
  wire [2:0] _T_88413; // @[AxiLoadQueue.scala 191:60:@35227.4]
  wire [2:0] _T_88414; // @[AxiLoadQueue.scala 191:60:@35228.4]
  wire [2:0] _T_88415; // @[AxiLoadQueue.scala 191:60:@35229.4]
  wire [3:0] _T_88416; // @[AxiLoadQueue.scala 191:60:@35230.4]
  wire [3:0] _T_88417; // @[AxiLoadQueue.scala 191:60:@35231.4]
  wire [3:0] _T_88418; // @[AxiLoadQueue.scala 191:60:@35232.4]
  wire [3:0] _T_88419; // @[AxiLoadQueue.scala 191:60:@35233.4]
  wire [3:0] _T_88420; // @[AxiLoadQueue.scala 191:60:@35234.4]
  wire [3:0] _T_88421; // @[AxiLoadQueue.scala 191:60:@35235.4]
  wire [3:0] _T_88422; // @[AxiLoadQueue.scala 191:60:@35236.4]
  wire [3:0] _T_88423; // @[AxiLoadQueue.scala 191:60:@35237.4]
  wire  _T_88426; // @[AxiLoadQueue.scala 192:43:@35239.4]
  wire  _T_88427; // @[AxiLoadQueue.scala 192:43:@35240.4]
  wire  _T_88428; // @[AxiLoadQueue.scala 192:43:@35241.4]
  wire  _T_88429; // @[AxiLoadQueue.scala 192:43:@35242.4]
  wire  _T_88430; // @[AxiLoadQueue.scala 192:43:@35243.4]
  wire  _T_88431; // @[AxiLoadQueue.scala 192:43:@35244.4]
  wire  _T_88432; // @[AxiLoadQueue.scala 192:43:@35245.4]
  wire  _T_88433; // @[AxiLoadQueue.scala 192:43:@35246.4]
  wire  _T_88434; // @[AxiLoadQueue.scala 192:43:@35247.4]
  wire  _T_88435; // @[AxiLoadQueue.scala 192:43:@35248.4]
  wire  _T_88436; // @[AxiLoadQueue.scala 192:43:@35249.4]
  wire  _T_88437; // @[AxiLoadQueue.scala 192:43:@35250.4]
  wire  _T_88438; // @[AxiLoadQueue.scala 192:43:@35251.4]
  wire  _T_88439; // @[AxiLoadQueue.scala 192:43:@35252.4]
  wire  _T_88440; // @[AxiLoadQueue.scala 192:43:@35253.4]
  wire  _GEN_930; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_931; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_932; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_933; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_934; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_935; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_936; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_937; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_938; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_939; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_940; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_941; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_942; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_943; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_944; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_945; // @[AxiLoadQueue.scala 193:43:@35255.6]
  wire  _GEN_947; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_948; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_949; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_950; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_951; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_952; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_953; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_954; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_955; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_956; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_957; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_958; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_959; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_960; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire  _GEN_961; // @[AxiLoadQueue.scala 194:31:@35256.6]
  wire [31:0] _GEN_963; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_964; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_965; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_966; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_967; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_968; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_969; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_970; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_971; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_972; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_973; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_974; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_975; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_976; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire [31:0] _GEN_977; // @[AxiLoadQueue.scala 195:31:@35257.6]
  wire  lastConflict_1_0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_1; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_2; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_3; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_4; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_5; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_6; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_7; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_8; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_9; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_10; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_11; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_12; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_13; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_14; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  lastConflict_1_15; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire  canBypass_1; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire [31:0] bypassVal_1; // @[AxiLoadQueue.scala 192:53:@35254.4]
  wire [1:0] _T_88546; // @[AxiLoadQueue.scala 191:60:@35311.4]
  wire [1:0] _T_88547; // @[AxiLoadQueue.scala 191:60:@35312.4]
  wire [2:0] _T_88548; // @[AxiLoadQueue.scala 191:60:@35313.4]
  wire [2:0] _T_88549; // @[AxiLoadQueue.scala 191:60:@35314.4]
  wire [2:0] _T_88550; // @[AxiLoadQueue.scala 191:60:@35315.4]
  wire [2:0] _T_88551; // @[AxiLoadQueue.scala 191:60:@35316.4]
  wire [3:0] _T_88552; // @[AxiLoadQueue.scala 191:60:@35317.4]
  wire [3:0] _T_88553; // @[AxiLoadQueue.scala 191:60:@35318.4]
  wire [3:0] _T_88554; // @[AxiLoadQueue.scala 191:60:@35319.4]
  wire [3:0] _T_88555; // @[AxiLoadQueue.scala 191:60:@35320.4]
  wire [3:0] _T_88556; // @[AxiLoadQueue.scala 191:60:@35321.4]
  wire [3:0] _T_88557; // @[AxiLoadQueue.scala 191:60:@35322.4]
  wire [3:0] _T_88558; // @[AxiLoadQueue.scala 191:60:@35323.4]
  wire [3:0] _T_88559; // @[AxiLoadQueue.scala 191:60:@35324.4]
  wire  _T_88562; // @[AxiLoadQueue.scala 192:43:@35326.4]
  wire  _T_88563; // @[AxiLoadQueue.scala 192:43:@35327.4]
  wire  _T_88564; // @[AxiLoadQueue.scala 192:43:@35328.4]
  wire  _T_88565; // @[AxiLoadQueue.scala 192:43:@35329.4]
  wire  _T_88566; // @[AxiLoadQueue.scala 192:43:@35330.4]
  wire  _T_88567; // @[AxiLoadQueue.scala 192:43:@35331.4]
  wire  _T_88568; // @[AxiLoadQueue.scala 192:43:@35332.4]
  wire  _T_88569; // @[AxiLoadQueue.scala 192:43:@35333.4]
  wire  _T_88570; // @[AxiLoadQueue.scala 192:43:@35334.4]
  wire  _T_88571; // @[AxiLoadQueue.scala 192:43:@35335.4]
  wire  _T_88572; // @[AxiLoadQueue.scala 192:43:@35336.4]
  wire  _T_88573; // @[AxiLoadQueue.scala 192:43:@35337.4]
  wire  _T_88574; // @[AxiLoadQueue.scala 192:43:@35338.4]
  wire  _T_88575; // @[AxiLoadQueue.scala 192:43:@35339.4]
  wire  _T_88576; // @[AxiLoadQueue.scala 192:43:@35340.4]
  wire  _GEN_996; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_997; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_998; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_999; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1000; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1001; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1002; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1003; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1004; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1005; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1006; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1007; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1008; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1009; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1010; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1011; // @[AxiLoadQueue.scala 193:43:@35342.6]
  wire  _GEN_1013; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1014; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1015; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1016; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1017; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1018; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1019; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1020; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1021; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1022; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1023; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1024; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1025; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1026; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire  _GEN_1027; // @[AxiLoadQueue.scala 194:31:@35343.6]
  wire [31:0] _GEN_1029; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1030; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1031; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1032; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1033; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1034; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1035; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1036; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1037; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1038; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1039; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1040; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1041; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1042; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire [31:0] _GEN_1043; // @[AxiLoadQueue.scala 195:31:@35344.6]
  wire  lastConflict_2_0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_1; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_2; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_3; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_4; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_5; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_6; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_7; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_8; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_9; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_10; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_11; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_12; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_13; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_14; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  lastConflict_2_15; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire  canBypass_2; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire [31:0] bypassVal_2; // @[AxiLoadQueue.scala 192:53:@35341.4]
  wire [1:0] _T_88682; // @[AxiLoadQueue.scala 191:60:@35398.4]
  wire [1:0] _T_88683; // @[AxiLoadQueue.scala 191:60:@35399.4]
  wire [2:0] _T_88684; // @[AxiLoadQueue.scala 191:60:@35400.4]
  wire [2:0] _T_88685; // @[AxiLoadQueue.scala 191:60:@35401.4]
  wire [2:0] _T_88686; // @[AxiLoadQueue.scala 191:60:@35402.4]
  wire [2:0] _T_88687; // @[AxiLoadQueue.scala 191:60:@35403.4]
  wire [3:0] _T_88688; // @[AxiLoadQueue.scala 191:60:@35404.4]
  wire [3:0] _T_88689; // @[AxiLoadQueue.scala 191:60:@35405.4]
  wire [3:0] _T_88690; // @[AxiLoadQueue.scala 191:60:@35406.4]
  wire [3:0] _T_88691; // @[AxiLoadQueue.scala 191:60:@35407.4]
  wire [3:0] _T_88692; // @[AxiLoadQueue.scala 191:60:@35408.4]
  wire [3:0] _T_88693; // @[AxiLoadQueue.scala 191:60:@35409.4]
  wire [3:0] _T_88694; // @[AxiLoadQueue.scala 191:60:@35410.4]
  wire [3:0] _T_88695; // @[AxiLoadQueue.scala 191:60:@35411.4]
  wire  _T_88698; // @[AxiLoadQueue.scala 192:43:@35413.4]
  wire  _T_88699; // @[AxiLoadQueue.scala 192:43:@35414.4]
  wire  _T_88700; // @[AxiLoadQueue.scala 192:43:@35415.4]
  wire  _T_88701; // @[AxiLoadQueue.scala 192:43:@35416.4]
  wire  _T_88702; // @[AxiLoadQueue.scala 192:43:@35417.4]
  wire  _T_88703; // @[AxiLoadQueue.scala 192:43:@35418.4]
  wire  _T_88704; // @[AxiLoadQueue.scala 192:43:@35419.4]
  wire  _T_88705; // @[AxiLoadQueue.scala 192:43:@35420.4]
  wire  _T_88706; // @[AxiLoadQueue.scala 192:43:@35421.4]
  wire  _T_88707; // @[AxiLoadQueue.scala 192:43:@35422.4]
  wire  _T_88708; // @[AxiLoadQueue.scala 192:43:@35423.4]
  wire  _T_88709; // @[AxiLoadQueue.scala 192:43:@35424.4]
  wire  _T_88710; // @[AxiLoadQueue.scala 192:43:@35425.4]
  wire  _T_88711; // @[AxiLoadQueue.scala 192:43:@35426.4]
  wire  _T_88712; // @[AxiLoadQueue.scala 192:43:@35427.4]
  wire  _GEN_1062; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1063; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1064; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1065; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1066; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1067; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1068; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1069; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1070; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1071; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1072; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1073; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1074; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1075; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1076; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1077; // @[AxiLoadQueue.scala 193:43:@35429.6]
  wire  _GEN_1079; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1080; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1081; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1082; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1083; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1084; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1085; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1086; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1087; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1088; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1089; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1090; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1091; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1092; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire  _GEN_1093; // @[AxiLoadQueue.scala 194:31:@35430.6]
  wire [31:0] _GEN_1095; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1096; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1097; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1098; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1099; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1100; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1101; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1102; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1103; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1104; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1105; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1106; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1107; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1108; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire [31:0] _GEN_1109; // @[AxiLoadQueue.scala 195:31:@35431.6]
  wire  lastConflict_3_0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_1; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_2; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_3; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_4; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_5; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_6; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_7; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_8; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_9; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_10; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_11; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_12; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_13; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_14; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  lastConflict_3_15; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire  canBypass_3; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire [31:0] bypassVal_3; // @[AxiLoadQueue.scala 192:53:@35428.4]
  wire [1:0] _T_88818; // @[AxiLoadQueue.scala 191:60:@35485.4]
  wire [1:0] _T_88819; // @[AxiLoadQueue.scala 191:60:@35486.4]
  wire [2:0] _T_88820; // @[AxiLoadQueue.scala 191:60:@35487.4]
  wire [2:0] _T_88821; // @[AxiLoadQueue.scala 191:60:@35488.4]
  wire [2:0] _T_88822; // @[AxiLoadQueue.scala 191:60:@35489.4]
  wire [2:0] _T_88823; // @[AxiLoadQueue.scala 191:60:@35490.4]
  wire [3:0] _T_88824; // @[AxiLoadQueue.scala 191:60:@35491.4]
  wire [3:0] _T_88825; // @[AxiLoadQueue.scala 191:60:@35492.4]
  wire [3:0] _T_88826; // @[AxiLoadQueue.scala 191:60:@35493.4]
  wire [3:0] _T_88827; // @[AxiLoadQueue.scala 191:60:@35494.4]
  wire [3:0] _T_88828; // @[AxiLoadQueue.scala 191:60:@35495.4]
  wire [3:0] _T_88829; // @[AxiLoadQueue.scala 191:60:@35496.4]
  wire [3:0] _T_88830; // @[AxiLoadQueue.scala 191:60:@35497.4]
  wire [3:0] _T_88831; // @[AxiLoadQueue.scala 191:60:@35498.4]
  wire  _T_88834; // @[AxiLoadQueue.scala 192:43:@35500.4]
  wire  _T_88835; // @[AxiLoadQueue.scala 192:43:@35501.4]
  wire  _T_88836; // @[AxiLoadQueue.scala 192:43:@35502.4]
  wire  _T_88837; // @[AxiLoadQueue.scala 192:43:@35503.4]
  wire  _T_88838; // @[AxiLoadQueue.scala 192:43:@35504.4]
  wire  _T_88839; // @[AxiLoadQueue.scala 192:43:@35505.4]
  wire  _T_88840; // @[AxiLoadQueue.scala 192:43:@35506.4]
  wire  _T_88841; // @[AxiLoadQueue.scala 192:43:@35507.4]
  wire  _T_88842; // @[AxiLoadQueue.scala 192:43:@35508.4]
  wire  _T_88843; // @[AxiLoadQueue.scala 192:43:@35509.4]
  wire  _T_88844; // @[AxiLoadQueue.scala 192:43:@35510.4]
  wire  _T_88845; // @[AxiLoadQueue.scala 192:43:@35511.4]
  wire  _T_88846; // @[AxiLoadQueue.scala 192:43:@35512.4]
  wire  _T_88847; // @[AxiLoadQueue.scala 192:43:@35513.4]
  wire  _T_88848; // @[AxiLoadQueue.scala 192:43:@35514.4]
  wire  _GEN_1128; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1129; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1130; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1131; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1132; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1133; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1134; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1135; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1136; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1137; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1138; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1139; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1140; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1141; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1142; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1143; // @[AxiLoadQueue.scala 193:43:@35516.6]
  wire  _GEN_1145; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1146; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1147; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1148; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1149; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1150; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1151; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1152; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1153; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1154; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1155; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1156; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1157; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1158; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire  _GEN_1159; // @[AxiLoadQueue.scala 194:31:@35517.6]
  wire [31:0] _GEN_1161; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1162; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1163; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1164; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1165; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1166; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1167; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1168; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1169; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1170; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1171; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1172; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1173; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1174; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire [31:0] _GEN_1175; // @[AxiLoadQueue.scala 195:31:@35518.6]
  wire  lastConflict_4_0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_1; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_2; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_3; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_4; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_5; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_6; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_7; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_8; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_9; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_10; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_11; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_12; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_13; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_14; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  lastConflict_4_15; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire  canBypass_4; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire [31:0] bypassVal_4; // @[AxiLoadQueue.scala 192:53:@35515.4]
  wire [1:0] _T_88954; // @[AxiLoadQueue.scala 191:60:@35572.4]
  wire [1:0] _T_88955; // @[AxiLoadQueue.scala 191:60:@35573.4]
  wire [2:0] _T_88956; // @[AxiLoadQueue.scala 191:60:@35574.4]
  wire [2:0] _T_88957; // @[AxiLoadQueue.scala 191:60:@35575.4]
  wire [2:0] _T_88958; // @[AxiLoadQueue.scala 191:60:@35576.4]
  wire [2:0] _T_88959; // @[AxiLoadQueue.scala 191:60:@35577.4]
  wire [3:0] _T_88960; // @[AxiLoadQueue.scala 191:60:@35578.4]
  wire [3:0] _T_88961; // @[AxiLoadQueue.scala 191:60:@35579.4]
  wire [3:0] _T_88962; // @[AxiLoadQueue.scala 191:60:@35580.4]
  wire [3:0] _T_88963; // @[AxiLoadQueue.scala 191:60:@35581.4]
  wire [3:0] _T_88964; // @[AxiLoadQueue.scala 191:60:@35582.4]
  wire [3:0] _T_88965; // @[AxiLoadQueue.scala 191:60:@35583.4]
  wire [3:0] _T_88966; // @[AxiLoadQueue.scala 191:60:@35584.4]
  wire [3:0] _T_88967; // @[AxiLoadQueue.scala 191:60:@35585.4]
  wire  _T_88970; // @[AxiLoadQueue.scala 192:43:@35587.4]
  wire  _T_88971; // @[AxiLoadQueue.scala 192:43:@35588.4]
  wire  _T_88972; // @[AxiLoadQueue.scala 192:43:@35589.4]
  wire  _T_88973; // @[AxiLoadQueue.scala 192:43:@35590.4]
  wire  _T_88974; // @[AxiLoadQueue.scala 192:43:@35591.4]
  wire  _T_88975; // @[AxiLoadQueue.scala 192:43:@35592.4]
  wire  _T_88976; // @[AxiLoadQueue.scala 192:43:@35593.4]
  wire  _T_88977; // @[AxiLoadQueue.scala 192:43:@35594.4]
  wire  _T_88978; // @[AxiLoadQueue.scala 192:43:@35595.4]
  wire  _T_88979; // @[AxiLoadQueue.scala 192:43:@35596.4]
  wire  _T_88980; // @[AxiLoadQueue.scala 192:43:@35597.4]
  wire  _T_88981; // @[AxiLoadQueue.scala 192:43:@35598.4]
  wire  _T_88982; // @[AxiLoadQueue.scala 192:43:@35599.4]
  wire  _T_88983; // @[AxiLoadQueue.scala 192:43:@35600.4]
  wire  _T_88984; // @[AxiLoadQueue.scala 192:43:@35601.4]
  wire  _GEN_1194; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1195; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1196; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1197; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1198; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1199; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1200; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1201; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1202; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1203; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1204; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1205; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1206; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1207; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1208; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1209; // @[AxiLoadQueue.scala 193:43:@35603.6]
  wire  _GEN_1211; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1212; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1213; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1214; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1215; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1216; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1217; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1218; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1219; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1220; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1221; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1222; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1223; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1224; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire  _GEN_1225; // @[AxiLoadQueue.scala 194:31:@35604.6]
  wire [31:0] _GEN_1227; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1228; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1229; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1230; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1231; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1232; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1233; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1234; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1235; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1236; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1237; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1238; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1239; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1240; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire [31:0] _GEN_1241; // @[AxiLoadQueue.scala 195:31:@35605.6]
  wire  lastConflict_5_0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_1; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_2; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_3; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_4; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_5; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_6; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_7; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_8; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_9; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_10; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_11; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_12; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_13; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_14; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  lastConflict_5_15; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire  canBypass_5; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire [31:0] bypassVal_5; // @[AxiLoadQueue.scala 192:53:@35602.4]
  wire [1:0] _T_89090; // @[AxiLoadQueue.scala 191:60:@35659.4]
  wire [1:0] _T_89091; // @[AxiLoadQueue.scala 191:60:@35660.4]
  wire [2:0] _T_89092; // @[AxiLoadQueue.scala 191:60:@35661.4]
  wire [2:0] _T_89093; // @[AxiLoadQueue.scala 191:60:@35662.4]
  wire [2:0] _T_89094; // @[AxiLoadQueue.scala 191:60:@35663.4]
  wire [2:0] _T_89095; // @[AxiLoadQueue.scala 191:60:@35664.4]
  wire [3:0] _T_89096; // @[AxiLoadQueue.scala 191:60:@35665.4]
  wire [3:0] _T_89097; // @[AxiLoadQueue.scala 191:60:@35666.4]
  wire [3:0] _T_89098; // @[AxiLoadQueue.scala 191:60:@35667.4]
  wire [3:0] _T_89099; // @[AxiLoadQueue.scala 191:60:@35668.4]
  wire [3:0] _T_89100; // @[AxiLoadQueue.scala 191:60:@35669.4]
  wire [3:0] _T_89101; // @[AxiLoadQueue.scala 191:60:@35670.4]
  wire [3:0] _T_89102; // @[AxiLoadQueue.scala 191:60:@35671.4]
  wire [3:0] _T_89103; // @[AxiLoadQueue.scala 191:60:@35672.4]
  wire  _T_89106; // @[AxiLoadQueue.scala 192:43:@35674.4]
  wire  _T_89107; // @[AxiLoadQueue.scala 192:43:@35675.4]
  wire  _T_89108; // @[AxiLoadQueue.scala 192:43:@35676.4]
  wire  _T_89109; // @[AxiLoadQueue.scala 192:43:@35677.4]
  wire  _T_89110; // @[AxiLoadQueue.scala 192:43:@35678.4]
  wire  _T_89111; // @[AxiLoadQueue.scala 192:43:@35679.4]
  wire  _T_89112; // @[AxiLoadQueue.scala 192:43:@35680.4]
  wire  _T_89113; // @[AxiLoadQueue.scala 192:43:@35681.4]
  wire  _T_89114; // @[AxiLoadQueue.scala 192:43:@35682.4]
  wire  _T_89115; // @[AxiLoadQueue.scala 192:43:@35683.4]
  wire  _T_89116; // @[AxiLoadQueue.scala 192:43:@35684.4]
  wire  _T_89117; // @[AxiLoadQueue.scala 192:43:@35685.4]
  wire  _T_89118; // @[AxiLoadQueue.scala 192:43:@35686.4]
  wire  _T_89119; // @[AxiLoadQueue.scala 192:43:@35687.4]
  wire  _T_89120; // @[AxiLoadQueue.scala 192:43:@35688.4]
  wire  _GEN_1260; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1261; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1262; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1263; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1264; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1265; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1266; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1267; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1268; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1269; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1270; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1271; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1272; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1273; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1274; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1275; // @[AxiLoadQueue.scala 193:43:@35690.6]
  wire  _GEN_1277; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1278; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1279; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1280; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1281; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1282; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1283; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1284; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1285; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1286; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1287; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1288; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1289; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1290; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire  _GEN_1291; // @[AxiLoadQueue.scala 194:31:@35691.6]
  wire [31:0] _GEN_1293; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1294; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1295; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1296; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1297; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1298; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1299; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1300; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1301; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1302; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1303; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1304; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1305; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1306; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire [31:0] _GEN_1307; // @[AxiLoadQueue.scala 195:31:@35692.6]
  wire  lastConflict_6_0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_1; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_2; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_3; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_4; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_5; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_6; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_7; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_8; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_9; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_10; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_11; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_12; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_13; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_14; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  lastConflict_6_15; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire  canBypass_6; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire [31:0] bypassVal_6; // @[AxiLoadQueue.scala 192:53:@35689.4]
  wire [1:0] _T_89226; // @[AxiLoadQueue.scala 191:60:@35746.4]
  wire [1:0] _T_89227; // @[AxiLoadQueue.scala 191:60:@35747.4]
  wire [2:0] _T_89228; // @[AxiLoadQueue.scala 191:60:@35748.4]
  wire [2:0] _T_89229; // @[AxiLoadQueue.scala 191:60:@35749.4]
  wire [2:0] _T_89230; // @[AxiLoadQueue.scala 191:60:@35750.4]
  wire [2:0] _T_89231; // @[AxiLoadQueue.scala 191:60:@35751.4]
  wire [3:0] _T_89232; // @[AxiLoadQueue.scala 191:60:@35752.4]
  wire [3:0] _T_89233; // @[AxiLoadQueue.scala 191:60:@35753.4]
  wire [3:0] _T_89234; // @[AxiLoadQueue.scala 191:60:@35754.4]
  wire [3:0] _T_89235; // @[AxiLoadQueue.scala 191:60:@35755.4]
  wire [3:0] _T_89236; // @[AxiLoadQueue.scala 191:60:@35756.4]
  wire [3:0] _T_89237; // @[AxiLoadQueue.scala 191:60:@35757.4]
  wire [3:0] _T_89238; // @[AxiLoadQueue.scala 191:60:@35758.4]
  wire [3:0] _T_89239; // @[AxiLoadQueue.scala 191:60:@35759.4]
  wire  _T_89242; // @[AxiLoadQueue.scala 192:43:@35761.4]
  wire  _T_89243; // @[AxiLoadQueue.scala 192:43:@35762.4]
  wire  _T_89244; // @[AxiLoadQueue.scala 192:43:@35763.4]
  wire  _T_89245; // @[AxiLoadQueue.scala 192:43:@35764.4]
  wire  _T_89246; // @[AxiLoadQueue.scala 192:43:@35765.4]
  wire  _T_89247; // @[AxiLoadQueue.scala 192:43:@35766.4]
  wire  _T_89248; // @[AxiLoadQueue.scala 192:43:@35767.4]
  wire  _T_89249; // @[AxiLoadQueue.scala 192:43:@35768.4]
  wire  _T_89250; // @[AxiLoadQueue.scala 192:43:@35769.4]
  wire  _T_89251; // @[AxiLoadQueue.scala 192:43:@35770.4]
  wire  _T_89252; // @[AxiLoadQueue.scala 192:43:@35771.4]
  wire  _T_89253; // @[AxiLoadQueue.scala 192:43:@35772.4]
  wire  _T_89254; // @[AxiLoadQueue.scala 192:43:@35773.4]
  wire  _T_89255; // @[AxiLoadQueue.scala 192:43:@35774.4]
  wire  _T_89256; // @[AxiLoadQueue.scala 192:43:@35775.4]
  wire  _GEN_1326; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1327; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1328; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1329; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1330; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1331; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1332; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1333; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1334; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1335; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1336; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1337; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1338; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1339; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1340; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1341; // @[AxiLoadQueue.scala 193:43:@35777.6]
  wire  _GEN_1343; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1344; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1345; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1346; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1347; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1348; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1349; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1350; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1351; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1352; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1353; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1354; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1355; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1356; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire  _GEN_1357; // @[AxiLoadQueue.scala 194:31:@35778.6]
  wire [31:0] _GEN_1359; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1360; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1361; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1362; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1363; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1364; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1365; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1366; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1367; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1368; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1369; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1370; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1371; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1372; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire [31:0] _GEN_1373; // @[AxiLoadQueue.scala 195:31:@35779.6]
  wire  lastConflict_7_0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_1; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_2; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_3; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_4; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_5; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_6; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_7; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_8; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_9; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_10; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_11; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_12; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_13; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_14; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  lastConflict_7_15; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire  canBypass_7; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire [31:0] bypassVal_7; // @[AxiLoadQueue.scala 192:53:@35776.4]
  wire [1:0] _T_89362; // @[AxiLoadQueue.scala 191:60:@35833.4]
  wire [1:0] _T_89363; // @[AxiLoadQueue.scala 191:60:@35834.4]
  wire [2:0] _T_89364; // @[AxiLoadQueue.scala 191:60:@35835.4]
  wire [2:0] _T_89365; // @[AxiLoadQueue.scala 191:60:@35836.4]
  wire [2:0] _T_89366; // @[AxiLoadQueue.scala 191:60:@35837.4]
  wire [2:0] _T_89367; // @[AxiLoadQueue.scala 191:60:@35838.4]
  wire [3:0] _T_89368; // @[AxiLoadQueue.scala 191:60:@35839.4]
  wire [3:0] _T_89369; // @[AxiLoadQueue.scala 191:60:@35840.4]
  wire [3:0] _T_89370; // @[AxiLoadQueue.scala 191:60:@35841.4]
  wire [3:0] _T_89371; // @[AxiLoadQueue.scala 191:60:@35842.4]
  wire [3:0] _T_89372; // @[AxiLoadQueue.scala 191:60:@35843.4]
  wire [3:0] _T_89373; // @[AxiLoadQueue.scala 191:60:@35844.4]
  wire [3:0] _T_89374; // @[AxiLoadQueue.scala 191:60:@35845.4]
  wire [3:0] _T_89375; // @[AxiLoadQueue.scala 191:60:@35846.4]
  wire  _T_89378; // @[AxiLoadQueue.scala 192:43:@35848.4]
  wire  _T_89379; // @[AxiLoadQueue.scala 192:43:@35849.4]
  wire  _T_89380; // @[AxiLoadQueue.scala 192:43:@35850.4]
  wire  _T_89381; // @[AxiLoadQueue.scala 192:43:@35851.4]
  wire  _T_89382; // @[AxiLoadQueue.scala 192:43:@35852.4]
  wire  _T_89383; // @[AxiLoadQueue.scala 192:43:@35853.4]
  wire  _T_89384; // @[AxiLoadQueue.scala 192:43:@35854.4]
  wire  _T_89385; // @[AxiLoadQueue.scala 192:43:@35855.4]
  wire  _T_89386; // @[AxiLoadQueue.scala 192:43:@35856.4]
  wire  _T_89387; // @[AxiLoadQueue.scala 192:43:@35857.4]
  wire  _T_89388; // @[AxiLoadQueue.scala 192:43:@35858.4]
  wire  _T_89389; // @[AxiLoadQueue.scala 192:43:@35859.4]
  wire  _T_89390; // @[AxiLoadQueue.scala 192:43:@35860.4]
  wire  _T_89391; // @[AxiLoadQueue.scala 192:43:@35861.4]
  wire  _T_89392; // @[AxiLoadQueue.scala 192:43:@35862.4]
  wire  _GEN_1392; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1393; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1394; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1395; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1396; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1397; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1398; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1399; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1400; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1401; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1402; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1403; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1404; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1405; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1406; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1407; // @[AxiLoadQueue.scala 193:43:@35864.6]
  wire  _GEN_1409; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1410; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1411; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1412; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1413; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1414; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1415; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1416; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1417; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1418; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1419; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1420; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1421; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1422; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire  _GEN_1423; // @[AxiLoadQueue.scala 194:31:@35865.6]
  wire [31:0] _GEN_1425; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1426; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1427; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1428; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1429; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1430; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1431; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1432; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1433; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1434; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1435; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1436; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1437; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1438; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire [31:0] _GEN_1439; // @[AxiLoadQueue.scala 195:31:@35866.6]
  wire  lastConflict_8_0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_1; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_2; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_3; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_4; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_5; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_6; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_7; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_8; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_9; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_10; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_11; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_12; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_13; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_14; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  lastConflict_8_15; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire  canBypass_8; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire [31:0] bypassVal_8; // @[AxiLoadQueue.scala 192:53:@35863.4]
  wire [1:0] _T_89498; // @[AxiLoadQueue.scala 191:60:@35920.4]
  wire [1:0] _T_89499; // @[AxiLoadQueue.scala 191:60:@35921.4]
  wire [2:0] _T_89500; // @[AxiLoadQueue.scala 191:60:@35922.4]
  wire [2:0] _T_89501; // @[AxiLoadQueue.scala 191:60:@35923.4]
  wire [2:0] _T_89502; // @[AxiLoadQueue.scala 191:60:@35924.4]
  wire [2:0] _T_89503; // @[AxiLoadQueue.scala 191:60:@35925.4]
  wire [3:0] _T_89504; // @[AxiLoadQueue.scala 191:60:@35926.4]
  wire [3:0] _T_89505; // @[AxiLoadQueue.scala 191:60:@35927.4]
  wire [3:0] _T_89506; // @[AxiLoadQueue.scala 191:60:@35928.4]
  wire [3:0] _T_89507; // @[AxiLoadQueue.scala 191:60:@35929.4]
  wire [3:0] _T_89508; // @[AxiLoadQueue.scala 191:60:@35930.4]
  wire [3:0] _T_89509; // @[AxiLoadQueue.scala 191:60:@35931.4]
  wire [3:0] _T_89510; // @[AxiLoadQueue.scala 191:60:@35932.4]
  wire [3:0] _T_89511; // @[AxiLoadQueue.scala 191:60:@35933.4]
  wire  _T_89514; // @[AxiLoadQueue.scala 192:43:@35935.4]
  wire  _T_89515; // @[AxiLoadQueue.scala 192:43:@35936.4]
  wire  _T_89516; // @[AxiLoadQueue.scala 192:43:@35937.4]
  wire  _T_89517; // @[AxiLoadQueue.scala 192:43:@35938.4]
  wire  _T_89518; // @[AxiLoadQueue.scala 192:43:@35939.4]
  wire  _T_89519; // @[AxiLoadQueue.scala 192:43:@35940.4]
  wire  _T_89520; // @[AxiLoadQueue.scala 192:43:@35941.4]
  wire  _T_89521; // @[AxiLoadQueue.scala 192:43:@35942.4]
  wire  _T_89522; // @[AxiLoadQueue.scala 192:43:@35943.4]
  wire  _T_89523; // @[AxiLoadQueue.scala 192:43:@35944.4]
  wire  _T_89524; // @[AxiLoadQueue.scala 192:43:@35945.4]
  wire  _T_89525; // @[AxiLoadQueue.scala 192:43:@35946.4]
  wire  _T_89526; // @[AxiLoadQueue.scala 192:43:@35947.4]
  wire  _T_89527; // @[AxiLoadQueue.scala 192:43:@35948.4]
  wire  _T_89528; // @[AxiLoadQueue.scala 192:43:@35949.4]
  wire  _GEN_1458; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1459; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1460; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1461; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1462; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1463; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1464; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1465; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1466; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1467; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1468; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1469; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1470; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1471; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1472; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1473; // @[AxiLoadQueue.scala 193:43:@35951.6]
  wire  _GEN_1475; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1476; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1477; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1478; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1479; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1480; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1481; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1482; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1483; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1484; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1485; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1486; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1487; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1488; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire  _GEN_1489; // @[AxiLoadQueue.scala 194:31:@35952.6]
  wire [31:0] _GEN_1491; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1492; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1493; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1494; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1495; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1496; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1497; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1498; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1499; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1500; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1501; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1502; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1503; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1504; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire [31:0] _GEN_1505; // @[AxiLoadQueue.scala 195:31:@35953.6]
  wire  lastConflict_9_0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_1; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_2; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_3; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_4; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_5; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_6; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_7; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_8; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_9; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_10; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_11; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_12; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_13; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_14; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  lastConflict_9_15; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire  canBypass_9; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire [31:0] bypassVal_9; // @[AxiLoadQueue.scala 192:53:@35950.4]
  wire [1:0] _T_89634; // @[AxiLoadQueue.scala 191:60:@36007.4]
  wire [1:0] _T_89635; // @[AxiLoadQueue.scala 191:60:@36008.4]
  wire [2:0] _T_89636; // @[AxiLoadQueue.scala 191:60:@36009.4]
  wire [2:0] _T_89637; // @[AxiLoadQueue.scala 191:60:@36010.4]
  wire [2:0] _T_89638; // @[AxiLoadQueue.scala 191:60:@36011.4]
  wire [2:0] _T_89639; // @[AxiLoadQueue.scala 191:60:@36012.4]
  wire [3:0] _T_89640; // @[AxiLoadQueue.scala 191:60:@36013.4]
  wire [3:0] _T_89641; // @[AxiLoadQueue.scala 191:60:@36014.4]
  wire [3:0] _T_89642; // @[AxiLoadQueue.scala 191:60:@36015.4]
  wire [3:0] _T_89643; // @[AxiLoadQueue.scala 191:60:@36016.4]
  wire [3:0] _T_89644; // @[AxiLoadQueue.scala 191:60:@36017.4]
  wire [3:0] _T_89645; // @[AxiLoadQueue.scala 191:60:@36018.4]
  wire [3:0] _T_89646; // @[AxiLoadQueue.scala 191:60:@36019.4]
  wire [3:0] _T_89647; // @[AxiLoadQueue.scala 191:60:@36020.4]
  wire  _T_89650; // @[AxiLoadQueue.scala 192:43:@36022.4]
  wire  _T_89651; // @[AxiLoadQueue.scala 192:43:@36023.4]
  wire  _T_89652; // @[AxiLoadQueue.scala 192:43:@36024.4]
  wire  _T_89653; // @[AxiLoadQueue.scala 192:43:@36025.4]
  wire  _T_89654; // @[AxiLoadQueue.scala 192:43:@36026.4]
  wire  _T_89655; // @[AxiLoadQueue.scala 192:43:@36027.4]
  wire  _T_89656; // @[AxiLoadQueue.scala 192:43:@36028.4]
  wire  _T_89657; // @[AxiLoadQueue.scala 192:43:@36029.4]
  wire  _T_89658; // @[AxiLoadQueue.scala 192:43:@36030.4]
  wire  _T_89659; // @[AxiLoadQueue.scala 192:43:@36031.4]
  wire  _T_89660; // @[AxiLoadQueue.scala 192:43:@36032.4]
  wire  _T_89661; // @[AxiLoadQueue.scala 192:43:@36033.4]
  wire  _T_89662; // @[AxiLoadQueue.scala 192:43:@36034.4]
  wire  _T_89663; // @[AxiLoadQueue.scala 192:43:@36035.4]
  wire  _T_89664; // @[AxiLoadQueue.scala 192:43:@36036.4]
  wire  _GEN_1524; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1525; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1526; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1527; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1528; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1529; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1530; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1531; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1532; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1533; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1534; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1535; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1536; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1537; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1538; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1539; // @[AxiLoadQueue.scala 193:43:@36038.6]
  wire  _GEN_1541; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1542; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1543; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1544; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1545; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1546; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1547; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1548; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1549; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1550; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1551; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1552; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1553; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1554; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire  _GEN_1555; // @[AxiLoadQueue.scala 194:31:@36039.6]
  wire [31:0] _GEN_1557; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1558; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1559; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1560; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1561; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1562; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1563; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1564; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1565; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1566; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1567; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1568; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1569; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1570; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire [31:0] _GEN_1571; // @[AxiLoadQueue.scala 195:31:@36040.6]
  wire  lastConflict_10_0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_1; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_2; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_3; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_4; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_5; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_6; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_7; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_8; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_9; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_10; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_11; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_12; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_13; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_14; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  lastConflict_10_15; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire  canBypass_10; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire [31:0] bypassVal_10; // @[AxiLoadQueue.scala 192:53:@36037.4]
  wire [1:0] _T_89770; // @[AxiLoadQueue.scala 191:60:@36094.4]
  wire [1:0] _T_89771; // @[AxiLoadQueue.scala 191:60:@36095.4]
  wire [2:0] _T_89772; // @[AxiLoadQueue.scala 191:60:@36096.4]
  wire [2:0] _T_89773; // @[AxiLoadQueue.scala 191:60:@36097.4]
  wire [2:0] _T_89774; // @[AxiLoadQueue.scala 191:60:@36098.4]
  wire [2:0] _T_89775; // @[AxiLoadQueue.scala 191:60:@36099.4]
  wire [3:0] _T_89776; // @[AxiLoadQueue.scala 191:60:@36100.4]
  wire [3:0] _T_89777; // @[AxiLoadQueue.scala 191:60:@36101.4]
  wire [3:0] _T_89778; // @[AxiLoadQueue.scala 191:60:@36102.4]
  wire [3:0] _T_89779; // @[AxiLoadQueue.scala 191:60:@36103.4]
  wire [3:0] _T_89780; // @[AxiLoadQueue.scala 191:60:@36104.4]
  wire [3:0] _T_89781; // @[AxiLoadQueue.scala 191:60:@36105.4]
  wire [3:0] _T_89782; // @[AxiLoadQueue.scala 191:60:@36106.4]
  wire [3:0] _T_89783; // @[AxiLoadQueue.scala 191:60:@36107.4]
  wire  _T_89786; // @[AxiLoadQueue.scala 192:43:@36109.4]
  wire  _T_89787; // @[AxiLoadQueue.scala 192:43:@36110.4]
  wire  _T_89788; // @[AxiLoadQueue.scala 192:43:@36111.4]
  wire  _T_89789; // @[AxiLoadQueue.scala 192:43:@36112.4]
  wire  _T_89790; // @[AxiLoadQueue.scala 192:43:@36113.4]
  wire  _T_89791; // @[AxiLoadQueue.scala 192:43:@36114.4]
  wire  _T_89792; // @[AxiLoadQueue.scala 192:43:@36115.4]
  wire  _T_89793; // @[AxiLoadQueue.scala 192:43:@36116.4]
  wire  _T_89794; // @[AxiLoadQueue.scala 192:43:@36117.4]
  wire  _T_89795; // @[AxiLoadQueue.scala 192:43:@36118.4]
  wire  _T_89796; // @[AxiLoadQueue.scala 192:43:@36119.4]
  wire  _T_89797; // @[AxiLoadQueue.scala 192:43:@36120.4]
  wire  _T_89798; // @[AxiLoadQueue.scala 192:43:@36121.4]
  wire  _T_89799; // @[AxiLoadQueue.scala 192:43:@36122.4]
  wire  _T_89800; // @[AxiLoadQueue.scala 192:43:@36123.4]
  wire  _GEN_1590; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1591; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1592; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1593; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1594; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1595; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1596; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1597; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1598; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1599; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1600; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1601; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1602; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1603; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1604; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1605; // @[AxiLoadQueue.scala 193:43:@36125.6]
  wire  _GEN_1607; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1608; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1609; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1610; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1611; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1612; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1613; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1614; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1615; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1616; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1617; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1618; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1619; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1620; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire  _GEN_1621; // @[AxiLoadQueue.scala 194:31:@36126.6]
  wire [31:0] _GEN_1623; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1624; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1625; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1626; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1627; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1628; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1629; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1630; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1631; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1632; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1633; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1634; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1635; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1636; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire [31:0] _GEN_1637; // @[AxiLoadQueue.scala 195:31:@36127.6]
  wire  lastConflict_11_0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_1; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_2; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_3; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_4; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_5; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_6; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_7; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_8; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_9; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_10; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_11; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_12; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_13; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_14; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  lastConflict_11_15; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire  canBypass_11; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire [31:0] bypassVal_11; // @[AxiLoadQueue.scala 192:53:@36124.4]
  wire [1:0] _T_89906; // @[AxiLoadQueue.scala 191:60:@36181.4]
  wire [1:0] _T_89907; // @[AxiLoadQueue.scala 191:60:@36182.4]
  wire [2:0] _T_89908; // @[AxiLoadQueue.scala 191:60:@36183.4]
  wire [2:0] _T_89909; // @[AxiLoadQueue.scala 191:60:@36184.4]
  wire [2:0] _T_89910; // @[AxiLoadQueue.scala 191:60:@36185.4]
  wire [2:0] _T_89911; // @[AxiLoadQueue.scala 191:60:@36186.4]
  wire [3:0] _T_89912; // @[AxiLoadQueue.scala 191:60:@36187.4]
  wire [3:0] _T_89913; // @[AxiLoadQueue.scala 191:60:@36188.4]
  wire [3:0] _T_89914; // @[AxiLoadQueue.scala 191:60:@36189.4]
  wire [3:0] _T_89915; // @[AxiLoadQueue.scala 191:60:@36190.4]
  wire [3:0] _T_89916; // @[AxiLoadQueue.scala 191:60:@36191.4]
  wire [3:0] _T_89917; // @[AxiLoadQueue.scala 191:60:@36192.4]
  wire [3:0] _T_89918; // @[AxiLoadQueue.scala 191:60:@36193.4]
  wire [3:0] _T_89919; // @[AxiLoadQueue.scala 191:60:@36194.4]
  wire  _T_89922; // @[AxiLoadQueue.scala 192:43:@36196.4]
  wire  _T_89923; // @[AxiLoadQueue.scala 192:43:@36197.4]
  wire  _T_89924; // @[AxiLoadQueue.scala 192:43:@36198.4]
  wire  _T_89925; // @[AxiLoadQueue.scala 192:43:@36199.4]
  wire  _T_89926; // @[AxiLoadQueue.scala 192:43:@36200.4]
  wire  _T_89927; // @[AxiLoadQueue.scala 192:43:@36201.4]
  wire  _T_89928; // @[AxiLoadQueue.scala 192:43:@36202.4]
  wire  _T_89929; // @[AxiLoadQueue.scala 192:43:@36203.4]
  wire  _T_89930; // @[AxiLoadQueue.scala 192:43:@36204.4]
  wire  _T_89931; // @[AxiLoadQueue.scala 192:43:@36205.4]
  wire  _T_89932; // @[AxiLoadQueue.scala 192:43:@36206.4]
  wire  _T_89933; // @[AxiLoadQueue.scala 192:43:@36207.4]
  wire  _T_89934; // @[AxiLoadQueue.scala 192:43:@36208.4]
  wire  _T_89935; // @[AxiLoadQueue.scala 192:43:@36209.4]
  wire  _T_89936; // @[AxiLoadQueue.scala 192:43:@36210.4]
  wire  _GEN_1656; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1657; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1658; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1659; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1660; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1661; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1662; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1663; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1664; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1665; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1666; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1667; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1668; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1669; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1670; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1671; // @[AxiLoadQueue.scala 193:43:@36212.6]
  wire  _GEN_1673; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1674; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1675; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1676; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1677; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1678; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1679; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1680; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1681; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1682; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1683; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1684; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1685; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1686; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire  _GEN_1687; // @[AxiLoadQueue.scala 194:31:@36213.6]
  wire [31:0] _GEN_1689; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1690; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1691; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1692; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1693; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1694; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1695; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1696; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1697; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1698; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1699; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1700; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1701; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1702; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire [31:0] _GEN_1703; // @[AxiLoadQueue.scala 195:31:@36214.6]
  wire  lastConflict_12_0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_1; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_2; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_3; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_4; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_5; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_6; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_7; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_8; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_9; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_10; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_11; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_12; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_13; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_14; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  lastConflict_12_15; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire  canBypass_12; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire [31:0] bypassVal_12; // @[AxiLoadQueue.scala 192:53:@36211.4]
  wire [1:0] _T_90042; // @[AxiLoadQueue.scala 191:60:@36268.4]
  wire [1:0] _T_90043; // @[AxiLoadQueue.scala 191:60:@36269.4]
  wire [2:0] _T_90044; // @[AxiLoadQueue.scala 191:60:@36270.4]
  wire [2:0] _T_90045; // @[AxiLoadQueue.scala 191:60:@36271.4]
  wire [2:0] _T_90046; // @[AxiLoadQueue.scala 191:60:@36272.4]
  wire [2:0] _T_90047; // @[AxiLoadQueue.scala 191:60:@36273.4]
  wire [3:0] _T_90048; // @[AxiLoadQueue.scala 191:60:@36274.4]
  wire [3:0] _T_90049; // @[AxiLoadQueue.scala 191:60:@36275.4]
  wire [3:0] _T_90050; // @[AxiLoadQueue.scala 191:60:@36276.4]
  wire [3:0] _T_90051; // @[AxiLoadQueue.scala 191:60:@36277.4]
  wire [3:0] _T_90052; // @[AxiLoadQueue.scala 191:60:@36278.4]
  wire [3:0] _T_90053; // @[AxiLoadQueue.scala 191:60:@36279.4]
  wire [3:0] _T_90054; // @[AxiLoadQueue.scala 191:60:@36280.4]
  wire [3:0] _T_90055; // @[AxiLoadQueue.scala 191:60:@36281.4]
  wire  _T_90058; // @[AxiLoadQueue.scala 192:43:@36283.4]
  wire  _T_90059; // @[AxiLoadQueue.scala 192:43:@36284.4]
  wire  _T_90060; // @[AxiLoadQueue.scala 192:43:@36285.4]
  wire  _T_90061; // @[AxiLoadQueue.scala 192:43:@36286.4]
  wire  _T_90062; // @[AxiLoadQueue.scala 192:43:@36287.4]
  wire  _T_90063; // @[AxiLoadQueue.scala 192:43:@36288.4]
  wire  _T_90064; // @[AxiLoadQueue.scala 192:43:@36289.4]
  wire  _T_90065; // @[AxiLoadQueue.scala 192:43:@36290.4]
  wire  _T_90066; // @[AxiLoadQueue.scala 192:43:@36291.4]
  wire  _T_90067; // @[AxiLoadQueue.scala 192:43:@36292.4]
  wire  _T_90068; // @[AxiLoadQueue.scala 192:43:@36293.4]
  wire  _T_90069; // @[AxiLoadQueue.scala 192:43:@36294.4]
  wire  _T_90070; // @[AxiLoadQueue.scala 192:43:@36295.4]
  wire  _T_90071; // @[AxiLoadQueue.scala 192:43:@36296.4]
  wire  _T_90072; // @[AxiLoadQueue.scala 192:43:@36297.4]
  wire  _GEN_1722; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1723; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1724; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1725; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1726; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1727; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1728; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1729; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1730; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1731; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1732; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1733; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1734; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1735; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1736; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1737; // @[AxiLoadQueue.scala 193:43:@36299.6]
  wire  _GEN_1739; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1740; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1741; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1742; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1743; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1744; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1745; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1746; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1747; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1748; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1749; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1750; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1751; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1752; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire  _GEN_1753; // @[AxiLoadQueue.scala 194:31:@36300.6]
  wire [31:0] _GEN_1755; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1756; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1757; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1758; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1759; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1760; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1761; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1762; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1763; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1764; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1765; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1766; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1767; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1768; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire [31:0] _GEN_1769; // @[AxiLoadQueue.scala 195:31:@36301.6]
  wire  lastConflict_13_0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_1; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_2; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_3; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_4; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_5; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_6; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_7; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_8; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_9; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_10; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_11; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_12; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_13; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_14; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  lastConflict_13_15; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire  canBypass_13; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire [31:0] bypassVal_13; // @[AxiLoadQueue.scala 192:53:@36298.4]
  wire [1:0] _T_90178; // @[AxiLoadQueue.scala 191:60:@36355.4]
  wire [1:0] _T_90179; // @[AxiLoadQueue.scala 191:60:@36356.4]
  wire [2:0] _T_90180; // @[AxiLoadQueue.scala 191:60:@36357.4]
  wire [2:0] _T_90181; // @[AxiLoadQueue.scala 191:60:@36358.4]
  wire [2:0] _T_90182; // @[AxiLoadQueue.scala 191:60:@36359.4]
  wire [2:0] _T_90183; // @[AxiLoadQueue.scala 191:60:@36360.4]
  wire [3:0] _T_90184; // @[AxiLoadQueue.scala 191:60:@36361.4]
  wire [3:0] _T_90185; // @[AxiLoadQueue.scala 191:60:@36362.4]
  wire [3:0] _T_90186; // @[AxiLoadQueue.scala 191:60:@36363.4]
  wire [3:0] _T_90187; // @[AxiLoadQueue.scala 191:60:@36364.4]
  wire [3:0] _T_90188; // @[AxiLoadQueue.scala 191:60:@36365.4]
  wire [3:0] _T_90189; // @[AxiLoadQueue.scala 191:60:@36366.4]
  wire [3:0] _T_90190; // @[AxiLoadQueue.scala 191:60:@36367.4]
  wire [3:0] _T_90191; // @[AxiLoadQueue.scala 191:60:@36368.4]
  wire  _T_90194; // @[AxiLoadQueue.scala 192:43:@36370.4]
  wire  _T_90195; // @[AxiLoadQueue.scala 192:43:@36371.4]
  wire  _T_90196; // @[AxiLoadQueue.scala 192:43:@36372.4]
  wire  _T_90197; // @[AxiLoadQueue.scala 192:43:@36373.4]
  wire  _T_90198; // @[AxiLoadQueue.scala 192:43:@36374.4]
  wire  _T_90199; // @[AxiLoadQueue.scala 192:43:@36375.4]
  wire  _T_90200; // @[AxiLoadQueue.scala 192:43:@36376.4]
  wire  _T_90201; // @[AxiLoadQueue.scala 192:43:@36377.4]
  wire  _T_90202; // @[AxiLoadQueue.scala 192:43:@36378.4]
  wire  _T_90203; // @[AxiLoadQueue.scala 192:43:@36379.4]
  wire  _T_90204; // @[AxiLoadQueue.scala 192:43:@36380.4]
  wire  _T_90205; // @[AxiLoadQueue.scala 192:43:@36381.4]
  wire  _T_90206; // @[AxiLoadQueue.scala 192:43:@36382.4]
  wire  _T_90207; // @[AxiLoadQueue.scala 192:43:@36383.4]
  wire  _T_90208; // @[AxiLoadQueue.scala 192:43:@36384.4]
  wire  _GEN_1788; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1789; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1790; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1791; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1792; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1793; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1794; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1795; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1796; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1797; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1798; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1799; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1800; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1801; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1802; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1803; // @[AxiLoadQueue.scala 193:43:@36386.6]
  wire  _GEN_1805; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1806; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1807; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1808; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1809; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1810; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1811; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1812; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1813; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1814; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1815; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1816; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1817; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1818; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire  _GEN_1819; // @[AxiLoadQueue.scala 194:31:@36387.6]
  wire [31:0] _GEN_1821; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1822; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1823; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1824; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1825; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1826; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1827; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1828; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1829; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1830; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1831; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1832; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1833; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1834; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire [31:0] _GEN_1835; // @[AxiLoadQueue.scala 195:31:@36388.6]
  wire  lastConflict_14_0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_1; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_2; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_3; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_4; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_5; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_6; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_7; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_8; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_9; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_10; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_11; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_12; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_13; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_14; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  lastConflict_14_15; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire  canBypass_14; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire [31:0] bypassVal_14; // @[AxiLoadQueue.scala 192:53:@36385.4]
  wire [1:0] _T_90314; // @[AxiLoadQueue.scala 191:60:@36442.4]
  wire [1:0] _T_90315; // @[AxiLoadQueue.scala 191:60:@36443.4]
  wire [2:0] _T_90316; // @[AxiLoadQueue.scala 191:60:@36444.4]
  wire [2:0] _T_90317; // @[AxiLoadQueue.scala 191:60:@36445.4]
  wire [2:0] _T_90318; // @[AxiLoadQueue.scala 191:60:@36446.4]
  wire [2:0] _T_90319; // @[AxiLoadQueue.scala 191:60:@36447.4]
  wire [3:0] _T_90320; // @[AxiLoadQueue.scala 191:60:@36448.4]
  wire [3:0] _T_90321; // @[AxiLoadQueue.scala 191:60:@36449.4]
  wire [3:0] _T_90322; // @[AxiLoadQueue.scala 191:60:@36450.4]
  wire [3:0] _T_90323; // @[AxiLoadQueue.scala 191:60:@36451.4]
  wire [3:0] _T_90324; // @[AxiLoadQueue.scala 191:60:@36452.4]
  wire [3:0] _T_90325; // @[AxiLoadQueue.scala 191:60:@36453.4]
  wire [3:0] _T_90326; // @[AxiLoadQueue.scala 191:60:@36454.4]
  wire [3:0] _T_90327; // @[AxiLoadQueue.scala 191:60:@36455.4]
  wire  _T_90330; // @[AxiLoadQueue.scala 192:43:@36457.4]
  wire  _T_90331; // @[AxiLoadQueue.scala 192:43:@36458.4]
  wire  _T_90332; // @[AxiLoadQueue.scala 192:43:@36459.4]
  wire  _T_90333; // @[AxiLoadQueue.scala 192:43:@36460.4]
  wire  _T_90334; // @[AxiLoadQueue.scala 192:43:@36461.4]
  wire  _T_90335; // @[AxiLoadQueue.scala 192:43:@36462.4]
  wire  _T_90336; // @[AxiLoadQueue.scala 192:43:@36463.4]
  wire  _T_90337; // @[AxiLoadQueue.scala 192:43:@36464.4]
  wire  _T_90338; // @[AxiLoadQueue.scala 192:43:@36465.4]
  wire  _T_90339; // @[AxiLoadQueue.scala 192:43:@36466.4]
  wire  _T_90340; // @[AxiLoadQueue.scala 192:43:@36467.4]
  wire  _T_90341; // @[AxiLoadQueue.scala 192:43:@36468.4]
  wire  _T_90342; // @[AxiLoadQueue.scala 192:43:@36469.4]
  wire  _T_90343; // @[AxiLoadQueue.scala 192:43:@36470.4]
  wire  _T_90344; // @[AxiLoadQueue.scala 192:43:@36471.4]
  wire  _GEN_1854; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1855; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1856; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1857; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1858; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1859; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1860; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1861; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1862; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1863; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1864; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1865; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1866; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1867; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1868; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1869; // @[AxiLoadQueue.scala 193:43:@36473.6]
  wire  _GEN_1871; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1872; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1873; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1874; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1875; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1876; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1877; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1878; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1879; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1880; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1881; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1882; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1883; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1884; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire  _GEN_1885; // @[AxiLoadQueue.scala 194:31:@36474.6]
  wire [31:0] _GEN_1887; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1888; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1889; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1890; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1891; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1892; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1893; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1894; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1895; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1896; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1897; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1898; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1899; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1900; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire [31:0] _GEN_1901; // @[AxiLoadQueue.scala 195:31:@36475.6]
  wire  lastConflict_15_0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_1; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_2; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_3; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_4; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_5; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_6; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_7; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_8; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_9; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_10; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_11; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_12; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_13; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_14; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  lastConflict_15_15; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire  canBypass_15; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire [31:0] bypassVal_15; // @[AxiLoadQueue.scala 192:53:@36472.4]
  wire [15:0] _T_90404; // @[OneHot.scala 52:12:@36480.4]
  wire  _T_90406; // @[util.scala 33:60:@36482.4]
  wire  _T_90407; // @[util.scala 33:60:@36483.4]
  wire  _T_90408; // @[util.scala 33:60:@36484.4]
  wire  _T_90409; // @[util.scala 33:60:@36485.4]
  wire  _T_90410; // @[util.scala 33:60:@36486.4]
  wire  _T_90411; // @[util.scala 33:60:@36487.4]
  wire  _T_90412; // @[util.scala 33:60:@36488.4]
  wire  _T_90413; // @[util.scala 33:60:@36489.4]
  wire  _T_90414; // @[util.scala 33:60:@36490.4]
  wire  _T_90415; // @[util.scala 33:60:@36491.4]
  wire  _T_90416; // @[util.scala 33:60:@36492.4]
  wire  _T_90417; // @[util.scala 33:60:@36493.4]
  wire  _T_90418; // @[util.scala 33:60:@36494.4]
  wire  _T_90419; // @[util.scala 33:60:@36495.4]
  wire  _T_90420; // @[util.scala 33:60:@36496.4]
  wire  _T_90421; // @[util.scala 33:60:@36497.4]
  wire  _T_93610; // @[AxiLoadQueue.scala 242:41:@39144.4]
  wire  _T_93611; // @[AxiLoadQueue.scala 242:38:@39145.4]
  wire  _T_93613; // @[AxiLoadQueue.scala 243:12:@39147.6]
  reg  loadInitiated_15; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_739;
  wire  _T_93615; // @[AxiLoadQueue.scala 243:46:@39148.6]
  wire  _T_93616; // @[AxiLoadQueue.scala 243:43:@39149.6]
  wire  _T_93618; // @[AxiLoadQueue.scala 243:78:@39150.6]
  wire  _T_93619; // @[AxiLoadQueue.scala 243:75:@39151.6]
  wire  _T_93622; // @[AxiLoadQueue.scala 246:86:@39154.8]
  wire  _T_93623; // @[AxiLoadQueue.scala 246:86:@39155.8]
  wire  _T_93624; // @[AxiLoadQueue.scala 246:86:@39156.8]
  wire  _T_93625; // @[AxiLoadQueue.scala 246:86:@39157.8]
  wire  _T_93626; // @[AxiLoadQueue.scala 246:86:@39158.8]
  wire  _T_93627; // @[AxiLoadQueue.scala 246:86:@39159.8]
  wire  _T_93628; // @[AxiLoadQueue.scala 246:86:@39160.8]
  wire  _T_93629; // @[AxiLoadQueue.scala 246:86:@39161.8]
  wire  _T_93630; // @[AxiLoadQueue.scala 246:86:@39162.8]
  wire  _T_93631; // @[AxiLoadQueue.scala 246:86:@39163.8]
  wire  _T_93632; // @[AxiLoadQueue.scala 246:86:@39164.8]
  wire  _T_93633; // @[AxiLoadQueue.scala 246:86:@39165.8]
  wire  _T_93634; // @[AxiLoadQueue.scala 246:86:@39166.8]
  wire  _T_93635; // @[AxiLoadQueue.scala 246:86:@39167.8]
  wire  _T_93636; // @[AxiLoadQueue.scala 246:86:@39168.8]
  wire  _T_93638; // @[AxiLoadQueue.scala 246:38:@39169.8]
  wire  _T_93657; // @[AxiLoadQueue.scala 247:11:@39186.8]
  wire  _T_93658; // @[AxiLoadQueue.scala 246:103:@39187.8]
  wire  _GEN_2060; // @[AxiLoadQueue.scala 243:104:@39152.6]
  wire  loadRequest_15; // @[AxiLoadQueue.scala 242:71:@39146.4]
  wire [15:0] _T_90462; // @[Mux.scala 31:69:@36515.4]
  wire  _T_93526; // @[AxiLoadQueue.scala 242:41:@39062.4]
  wire  _T_93527; // @[AxiLoadQueue.scala 242:38:@39063.4]
  wire  _T_93529; // @[AxiLoadQueue.scala 243:12:@39065.6]
  reg  loadInitiated_14; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_740;
  wire  _T_93531; // @[AxiLoadQueue.scala 243:46:@39066.6]
  wire  _T_93532; // @[AxiLoadQueue.scala 243:43:@39067.6]
  wire  _T_93534; // @[AxiLoadQueue.scala 243:78:@39068.6]
  wire  _T_93535; // @[AxiLoadQueue.scala 243:75:@39069.6]
  wire  _T_93538; // @[AxiLoadQueue.scala 246:86:@39072.8]
  wire  _T_93539; // @[AxiLoadQueue.scala 246:86:@39073.8]
  wire  _T_93540; // @[AxiLoadQueue.scala 246:86:@39074.8]
  wire  _T_93541; // @[AxiLoadQueue.scala 246:86:@39075.8]
  wire  _T_93542; // @[AxiLoadQueue.scala 246:86:@39076.8]
  wire  _T_93543; // @[AxiLoadQueue.scala 246:86:@39077.8]
  wire  _T_93544; // @[AxiLoadQueue.scala 246:86:@39078.8]
  wire  _T_93545; // @[AxiLoadQueue.scala 246:86:@39079.8]
  wire  _T_93546; // @[AxiLoadQueue.scala 246:86:@39080.8]
  wire  _T_93547; // @[AxiLoadQueue.scala 246:86:@39081.8]
  wire  _T_93548; // @[AxiLoadQueue.scala 246:86:@39082.8]
  wire  _T_93549; // @[AxiLoadQueue.scala 246:86:@39083.8]
  wire  _T_93550; // @[AxiLoadQueue.scala 246:86:@39084.8]
  wire  _T_93551; // @[AxiLoadQueue.scala 246:86:@39085.8]
  wire  _T_93552; // @[AxiLoadQueue.scala 246:86:@39086.8]
  wire  _T_93554; // @[AxiLoadQueue.scala 246:38:@39087.8]
  wire  _T_93573; // @[AxiLoadQueue.scala 247:11:@39104.8]
  wire  _T_93574; // @[AxiLoadQueue.scala 246:103:@39105.8]
  wire  _GEN_2056; // @[AxiLoadQueue.scala 243:104:@39070.6]
  wire  loadRequest_14; // @[AxiLoadQueue.scala 242:71:@39064.4]
  wire [15:0] _T_90463; // @[Mux.scala 31:69:@36516.4]
  wire  _T_93442; // @[AxiLoadQueue.scala 242:41:@38980.4]
  wire  _T_93443; // @[AxiLoadQueue.scala 242:38:@38981.4]
  wire  _T_93445; // @[AxiLoadQueue.scala 243:12:@38983.6]
  reg  loadInitiated_13; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_741;
  wire  _T_93447; // @[AxiLoadQueue.scala 243:46:@38984.6]
  wire  _T_93448; // @[AxiLoadQueue.scala 243:43:@38985.6]
  wire  _T_93450; // @[AxiLoadQueue.scala 243:78:@38986.6]
  wire  _T_93451; // @[AxiLoadQueue.scala 243:75:@38987.6]
  wire  _T_93454; // @[AxiLoadQueue.scala 246:86:@38990.8]
  wire  _T_93455; // @[AxiLoadQueue.scala 246:86:@38991.8]
  wire  _T_93456; // @[AxiLoadQueue.scala 246:86:@38992.8]
  wire  _T_93457; // @[AxiLoadQueue.scala 246:86:@38993.8]
  wire  _T_93458; // @[AxiLoadQueue.scala 246:86:@38994.8]
  wire  _T_93459; // @[AxiLoadQueue.scala 246:86:@38995.8]
  wire  _T_93460; // @[AxiLoadQueue.scala 246:86:@38996.8]
  wire  _T_93461; // @[AxiLoadQueue.scala 246:86:@38997.8]
  wire  _T_93462; // @[AxiLoadQueue.scala 246:86:@38998.8]
  wire  _T_93463; // @[AxiLoadQueue.scala 246:86:@38999.8]
  wire  _T_93464; // @[AxiLoadQueue.scala 246:86:@39000.8]
  wire  _T_93465; // @[AxiLoadQueue.scala 246:86:@39001.8]
  wire  _T_93466; // @[AxiLoadQueue.scala 246:86:@39002.8]
  wire  _T_93467; // @[AxiLoadQueue.scala 246:86:@39003.8]
  wire  _T_93468; // @[AxiLoadQueue.scala 246:86:@39004.8]
  wire  _T_93470; // @[AxiLoadQueue.scala 246:38:@39005.8]
  wire  _T_93489; // @[AxiLoadQueue.scala 247:11:@39022.8]
  wire  _T_93490; // @[AxiLoadQueue.scala 246:103:@39023.8]
  wire  _GEN_2052; // @[AxiLoadQueue.scala 243:104:@38988.6]
  wire  loadRequest_13; // @[AxiLoadQueue.scala 242:71:@38982.4]
  wire [15:0] _T_90464; // @[Mux.scala 31:69:@36517.4]
  wire  _T_93358; // @[AxiLoadQueue.scala 242:41:@38898.4]
  wire  _T_93359; // @[AxiLoadQueue.scala 242:38:@38899.4]
  wire  _T_93361; // @[AxiLoadQueue.scala 243:12:@38901.6]
  reg  loadInitiated_12; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_742;
  wire  _T_93363; // @[AxiLoadQueue.scala 243:46:@38902.6]
  wire  _T_93364; // @[AxiLoadQueue.scala 243:43:@38903.6]
  wire  _T_93366; // @[AxiLoadQueue.scala 243:78:@38904.6]
  wire  _T_93367; // @[AxiLoadQueue.scala 243:75:@38905.6]
  wire  _T_93370; // @[AxiLoadQueue.scala 246:86:@38908.8]
  wire  _T_93371; // @[AxiLoadQueue.scala 246:86:@38909.8]
  wire  _T_93372; // @[AxiLoadQueue.scala 246:86:@38910.8]
  wire  _T_93373; // @[AxiLoadQueue.scala 246:86:@38911.8]
  wire  _T_93374; // @[AxiLoadQueue.scala 246:86:@38912.8]
  wire  _T_93375; // @[AxiLoadQueue.scala 246:86:@38913.8]
  wire  _T_93376; // @[AxiLoadQueue.scala 246:86:@38914.8]
  wire  _T_93377; // @[AxiLoadQueue.scala 246:86:@38915.8]
  wire  _T_93378; // @[AxiLoadQueue.scala 246:86:@38916.8]
  wire  _T_93379; // @[AxiLoadQueue.scala 246:86:@38917.8]
  wire  _T_93380; // @[AxiLoadQueue.scala 246:86:@38918.8]
  wire  _T_93381; // @[AxiLoadQueue.scala 246:86:@38919.8]
  wire  _T_93382; // @[AxiLoadQueue.scala 246:86:@38920.8]
  wire  _T_93383; // @[AxiLoadQueue.scala 246:86:@38921.8]
  wire  _T_93384; // @[AxiLoadQueue.scala 246:86:@38922.8]
  wire  _T_93386; // @[AxiLoadQueue.scala 246:38:@38923.8]
  wire  _T_93405; // @[AxiLoadQueue.scala 247:11:@38940.8]
  wire  _T_93406; // @[AxiLoadQueue.scala 246:103:@38941.8]
  wire  _GEN_2048; // @[AxiLoadQueue.scala 243:104:@38906.6]
  wire  loadRequest_12; // @[AxiLoadQueue.scala 242:71:@38900.4]
  wire [15:0] _T_90465; // @[Mux.scala 31:69:@36518.4]
  wire  _T_93274; // @[AxiLoadQueue.scala 242:41:@38816.4]
  wire  _T_93275; // @[AxiLoadQueue.scala 242:38:@38817.4]
  wire  _T_93277; // @[AxiLoadQueue.scala 243:12:@38819.6]
  reg  loadInitiated_11; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_743;
  wire  _T_93279; // @[AxiLoadQueue.scala 243:46:@38820.6]
  wire  _T_93280; // @[AxiLoadQueue.scala 243:43:@38821.6]
  wire  _T_93282; // @[AxiLoadQueue.scala 243:78:@38822.6]
  wire  _T_93283; // @[AxiLoadQueue.scala 243:75:@38823.6]
  wire  _T_93286; // @[AxiLoadQueue.scala 246:86:@38826.8]
  wire  _T_93287; // @[AxiLoadQueue.scala 246:86:@38827.8]
  wire  _T_93288; // @[AxiLoadQueue.scala 246:86:@38828.8]
  wire  _T_93289; // @[AxiLoadQueue.scala 246:86:@38829.8]
  wire  _T_93290; // @[AxiLoadQueue.scala 246:86:@38830.8]
  wire  _T_93291; // @[AxiLoadQueue.scala 246:86:@38831.8]
  wire  _T_93292; // @[AxiLoadQueue.scala 246:86:@38832.8]
  wire  _T_93293; // @[AxiLoadQueue.scala 246:86:@38833.8]
  wire  _T_93294; // @[AxiLoadQueue.scala 246:86:@38834.8]
  wire  _T_93295; // @[AxiLoadQueue.scala 246:86:@38835.8]
  wire  _T_93296; // @[AxiLoadQueue.scala 246:86:@38836.8]
  wire  _T_93297; // @[AxiLoadQueue.scala 246:86:@38837.8]
  wire  _T_93298; // @[AxiLoadQueue.scala 246:86:@38838.8]
  wire  _T_93299; // @[AxiLoadQueue.scala 246:86:@38839.8]
  wire  _T_93300; // @[AxiLoadQueue.scala 246:86:@38840.8]
  wire  _T_93302; // @[AxiLoadQueue.scala 246:38:@38841.8]
  wire  _T_93321; // @[AxiLoadQueue.scala 247:11:@38858.8]
  wire  _T_93322; // @[AxiLoadQueue.scala 246:103:@38859.8]
  wire  _GEN_2044; // @[AxiLoadQueue.scala 243:104:@38824.6]
  wire  loadRequest_11; // @[AxiLoadQueue.scala 242:71:@38818.4]
  wire [15:0] _T_90466; // @[Mux.scala 31:69:@36519.4]
  wire  _T_93190; // @[AxiLoadQueue.scala 242:41:@38734.4]
  wire  _T_93191; // @[AxiLoadQueue.scala 242:38:@38735.4]
  wire  _T_93193; // @[AxiLoadQueue.scala 243:12:@38737.6]
  reg  loadInitiated_10; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_744;
  wire  _T_93195; // @[AxiLoadQueue.scala 243:46:@38738.6]
  wire  _T_93196; // @[AxiLoadQueue.scala 243:43:@38739.6]
  wire  _T_93198; // @[AxiLoadQueue.scala 243:78:@38740.6]
  wire  _T_93199; // @[AxiLoadQueue.scala 243:75:@38741.6]
  wire  _T_93202; // @[AxiLoadQueue.scala 246:86:@38744.8]
  wire  _T_93203; // @[AxiLoadQueue.scala 246:86:@38745.8]
  wire  _T_93204; // @[AxiLoadQueue.scala 246:86:@38746.8]
  wire  _T_93205; // @[AxiLoadQueue.scala 246:86:@38747.8]
  wire  _T_93206; // @[AxiLoadQueue.scala 246:86:@38748.8]
  wire  _T_93207; // @[AxiLoadQueue.scala 246:86:@38749.8]
  wire  _T_93208; // @[AxiLoadQueue.scala 246:86:@38750.8]
  wire  _T_93209; // @[AxiLoadQueue.scala 246:86:@38751.8]
  wire  _T_93210; // @[AxiLoadQueue.scala 246:86:@38752.8]
  wire  _T_93211; // @[AxiLoadQueue.scala 246:86:@38753.8]
  wire  _T_93212; // @[AxiLoadQueue.scala 246:86:@38754.8]
  wire  _T_93213; // @[AxiLoadQueue.scala 246:86:@38755.8]
  wire  _T_93214; // @[AxiLoadQueue.scala 246:86:@38756.8]
  wire  _T_93215; // @[AxiLoadQueue.scala 246:86:@38757.8]
  wire  _T_93216; // @[AxiLoadQueue.scala 246:86:@38758.8]
  wire  _T_93218; // @[AxiLoadQueue.scala 246:38:@38759.8]
  wire  _T_93237; // @[AxiLoadQueue.scala 247:11:@38776.8]
  wire  _T_93238; // @[AxiLoadQueue.scala 246:103:@38777.8]
  wire  _GEN_2040; // @[AxiLoadQueue.scala 243:104:@38742.6]
  wire  loadRequest_10; // @[AxiLoadQueue.scala 242:71:@38736.4]
  wire [15:0] _T_90467; // @[Mux.scala 31:69:@36520.4]
  wire  _T_93106; // @[AxiLoadQueue.scala 242:41:@38652.4]
  wire  _T_93107; // @[AxiLoadQueue.scala 242:38:@38653.4]
  wire  _T_93109; // @[AxiLoadQueue.scala 243:12:@38655.6]
  reg  loadInitiated_9; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_745;
  wire  _T_93111; // @[AxiLoadQueue.scala 243:46:@38656.6]
  wire  _T_93112; // @[AxiLoadQueue.scala 243:43:@38657.6]
  wire  _T_93114; // @[AxiLoadQueue.scala 243:78:@38658.6]
  wire  _T_93115; // @[AxiLoadQueue.scala 243:75:@38659.6]
  wire  _T_93118; // @[AxiLoadQueue.scala 246:86:@38662.8]
  wire  _T_93119; // @[AxiLoadQueue.scala 246:86:@38663.8]
  wire  _T_93120; // @[AxiLoadQueue.scala 246:86:@38664.8]
  wire  _T_93121; // @[AxiLoadQueue.scala 246:86:@38665.8]
  wire  _T_93122; // @[AxiLoadQueue.scala 246:86:@38666.8]
  wire  _T_93123; // @[AxiLoadQueue.scala 246:86:@38667.8]
  wire  _T_93124; // @[AxiLoadQueue.scala 246:86:@38668.8]
  wire  _T_93125; // @[AxiLoadQueue.scala 246:86:@38669.8]
  wire  _T_93126; // @[AxiLoadQueue.scala 246:86:@38670.8]
  wire  _T_93127; // @[AxiLoadQueue.scala 246:86:@38671.8]
  wire  _T_93128; // @[AxiLoadQueue.scala 246:86:@38672.8]
  wire  _T_93129; // @[AxiLoadQueue.scala 246:86:@38673.8]
  wire  _T_93130; // @[AxiLoadQueue.scala 246:86:@38674.8]
  wire  _T_93131; // @[AxiLoadQueue.scala 246:86:@38675.8]
  wire  _T_93132; // @[AxiLoadQueue.scala 246:86:@38676.8]
  wire  _T_93134; // @[AxiLoadQueue.scala 246:38:@38677.8]
  wire  _T_93153; // @[AxiLoadQueue.scala 247:11:@38694.8]
  wire  _T_93154; // @[AxiLoadQueue.scala 246:103:@38695.8]
  wire  _GEN_2036; // @[AxiLoadQueue.scala 243:104:@38660.6]
  wire  loadRequest_9; // @[AxiLoadQueue.scala 242:71:@38654.4]
  wire [15:0] _T_90468; // @[Mux.scala 31:69:@36521.4]
  wire  _T_93022; // @[AxiLoadQueue.scala 242:41:@38570.4]
  wire  _T_93023; // @[AxiLoadQueue.scala 242:38:@38571.4]
  wire  _T_93025; // @[AxiLoadQueue.scala 243:12:@38573.6]
  reg  loadInitiated_8; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_746;
  wire  _T_93027; // @[AxiLoadQueue.scala 243:46:@38574.6]
  wire  _T_93028; // @[AxiLoadQueue.scala 243:43:@38575.6]
  wire  _T_93030; // @[AxiLoadQueue.scala 243:78:@38576.6]
  wire  _T_93031; // @[AxiLoadQueue.scala 243:75:@38577.6]
  wire  _T_93034; // @[AxiLoadQueue.scala 246:86:@38580.8]
  wire  _T_93035; // @[AxiLoadQueue.scala 246:86:@38581.8]
  wire  _T_93036; // @[AxiLoadQueue.scala 246:86:@38582.8]
  wire  _T_93037; // @[AxiLoadQueue.scala 246:86:@38583.8]
  wire  _T_93038; // @[AxiLoadQueue.scala 246:86:@38584.8]
  wire  _T_93039; // @[AxiLoadQueue.scala 246:86:@38585.8]
  wire  _T_93040; // @[AxiLoadQueue.scala 246:86:@38586.8]
  wire  _T_93041; // @[AxiLoadQueue.scala 246:86:@38587.8]
  wire  _T_93042; // @[AxiLoadQueue.scala 246:86:@38588.8]
  wire  _T_93043; // @[AxiLoadQueue.scala 246:86:@38589.8]
  wire  _T_93044; // @[AxiLoadQueue.scala 246:86:@38590.8]
  wire  _T_93045; // @[AxiLoadQueue.scala 246:86:@38591.8]
  wire  _T_93046; // @[AxiLoadQueue.scala 246:86:@38592.8]
  wire  _T_93047; // @[AxiLoadQueue.scala 246:86:@38593.8]
  wire  _T_93048; // @[AxiLoadQueue.scala 246:86:@38594.8]
  wire  _T_93050; // @[AxiLoadQueue.scala 246:38:@38595.8]
  wire  _T_93069; // @[AxiLoadQueue.scala 247:11:@38612.8]
  wire  _T_93070; // @[AxiLoadQueue.scala 246:103:@38613.8]
  wire  _GEN_2032; // @[AxiLoadQueue.scala 243:104:@38578.6]
  wire  loadRequest_8; // @[AxiLoadQueue.scala 242:71:@38572.4]
  wire [15:0] _T_90469; // @[Mux.scala 31:69:@36522.4]
  wire  _T_92938; // @[AxiLoadQueue.scala 242:41:@38488.4]
  wire  _T_92939; // @[AxiLoadQueue.scala 242:38:@38489.4]
  wire  _T_92941; // @[AxiLoadQueue.scala 243:12:@38491.6]
  reg  loadInitiated_7; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_747;
  wire  _T_92943; // @[AxiLoadQueue.scala 243:46:@38492.6]
  wire  _T_92944; // @[AxiLoadQueue.scala 243:43:@38493.6]
  wire  _T_92946; // @[AxiLoadQueue.scala 243:78:@38494.6]
  wire  _T_92947; // @[AxiLoadQueue.scala 243:75:@38495.6]
  wire  _T_92950; // @[AxiLoadQueue.scala 246:86:@38498.8]
  wire  _T_92951; // @[AxiLoadQueue.scala 246:86:@38499.8]
  wire  _T_92952; // @[AxiLoadQueue.scala 246:86:@38500.8]
  wire  _T_92953; // @[AxiLoadQueue.scala 246:86:@38501.8]
  wire  _T_92954; // @[AxiLoadQueue.scala 246:86:@38502.8]
  wire  _T_92955; // @[AxiLoadQueue.scala 246:86:@38503.8]
  wire  _T_92956; // @[AxiLoadQueue.scala 246:86:@38504.8]
  wire  _T_92957; // @[AxiLoadQueue.scala 246:86:@38505.8]
  wire  _T_92958; // @[AxiLoadQueue.scala 246:86:@38506.8]
  wire  _T_92959; // @[AxiLoadQueue.scala 246:86:@38507.8]
  wire  _T_92960; // @[AxiLoadQueue.scala 246:86:@38508.8]
  wire  _T_92961; // @[AxiLoadQueue.scala 246:86:@38509.8]
  wire  _T_92962; // @[AxiLoadQueue.scala 246:86:@38510.8]
  wire  _T_92963; // @[AxiLoadQueue.scala 246:86:@38511.8]
  wire  _T_92964; // @[AxiLoadQueue.scala 246:86:@38512.8]
  wire  _T_92966; // @[AxiLoadQueue.scala 246:38:@38513.8]
  wire  _T_92985; // @[AxiLoadQueue.scala 247:11:@38530.8]
  wire  _T_92986; // @[AxiLoadQueue.scala 246:103:@38531.8]
  wire  _GEN_2028; // @[AxiLoadQueue.scala 243:104:@38496.6]
  wire  loadRequest_7; // @[AxiLoadQueue.scala 242:71:@38490.4]
  wire [15:0] _T_90470; // @[Mux.scala 31:69:@36523.4]
  wire  _T_92854; // @[AxiLoadQueue.scala 242:41:@38406.4]
  wire  _T_92855; // @[AxiLoadQueue.scala 242:38:@38407.4]
  wire  _T_92857; // @[AxiLoadQueue.scala 243:12:@38409.6]
  reg  loadInitiated_6; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_748;
  wire  _T_92859; // @[AxiLoadQueue.scala 243:46:@38410.6]
  wire  _T_92860; // @[AxiLoadQueue.scala 243:43:@38411.6]
  wire  _T_92862; // @[AxiLoadQueue.scala 243:78:@38412.6]
  wire  _T_92863; // @[AxiLoadQueue.scala 243:75:@38413.6]
  wire  _T_92866; // @[AxiLoadQueue.scala 246:86:@38416.8]
  wire  _T_92867; // @[AxiLoadQueue.scala 246:86:@38417.8]
  wire  _T_92868; // @[AxiLoadQueue.scala 246:86:@38418.8]
  wire  _T_92869; // @[AxiLoadQueue.scala 246:86:@38419.8]
  wire  _T_92870; // @[AxiLoadQueue.scala 246:86:@38420.8]
  wire  _T_92871; // @[AxiLoadQueue.scala 246:86:@38421.8]
  wire  _T_92872; // @[AxiLoadQueue.scala 246:86:@38422.8]
  wire  _T_92873; // @[AxiLoadQueue.scala 246:86:@38423.8]
  wire  _T_92874; // @[AxiLoadQueue.scala 246:86:@38424.8]
  wire  _T_92875; // @[AxiLoadQueue.scala 246:86:@38425.8]
  wire  _T_92876; // @[AxiLoadQueue.scala 246:86:@38426.8]
  wire  _T_92877; // @[AxiLoadQueue.scala 246:86:@38427.8]
  wire  _T_92878; // @[AxiLoadQueue.scala 246:86:@38428.8]
  wire  _T_92879; // @[AxiLoadQueue.scala 246:86:@38429.8]
  wire  _T_92880; // @[AxiLoadQueue.scala 246:86:@38430.8]
  wire  _T_92882; // @[AxiLoadQueue.scala 246:38:@38431.8]
  wire  _T_92901; // @[AxiLoadQueue.scala 247:11:@38448.8]
  wire  _T_92902; // @[AxiLoadQueue.scala 246:103:@38449.8]
  wire  _GEN_2024; // @[AxiLoadQueue.scala 243:104:@38414.6]
  wire  loadRequest_6; // @[AxiLoadQueue.scala 242:71:@38408.4]
  wire [15:0] _T_90471; // @[Mux.scala 31:69:@36524.4]
  wire  _T_92770; // @[AxiLoadQueue.scala 242:41:@38324.4]
  wire  _T_92771; // @[AxiLoadQueue.scala 242:38:@38325.4]
  wire  _T_92773; // @[AxiLoadQueue.scala 243:12:@38327.6]
  reg  loadInitiated_5; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_749;
  wire  _T_92775; // @[AxiLoadQueue.scala 243:46:@38328.6]
  wire  _T_92776; // @[AxiLoadQueue.scala 243:43:@38329.6]
  wire  _T_92778; // @[AxiLoadQueue.scala 243:78:@38330.6]
  wire  _T_92779; // @[AxiLoadQueue.scala 243:75:@38331.6]
  wire  _T_92782; // @[AxiLoadQueue.scala 246:86:@38334.8]
  wire  _T_92783; // @[AxiLoadQueue.scala 246:86:@38335.8]
  wire  _T_92784; // @[AxiLoadQueue.scala 246:86:@38336.8]
  wire  _T_92785; // @[AxiLoadQueue.scala 246:86:@38337.8]
  wire  _T_92786; // @[AxiLoadQueue.scala 246:86:@38338.8]
  wire  _T_92787; // @[AxiLoadQueue.scala 246:86:@38339.8]
  wire  _T_92788; // @[AxiLoadQueue.scala 246:86:@38340.8]
  wire  _T_92789; // @[AxiLoadQueue.scala 246:86:@38341.8]
  wire  _T_92790; // @[AxiLoadQueue.scala 246:86:@38342.8]
  wire  _T_92791; // @[AxiLoadQueue.scala 246:86:@38343.8]
  wire  _T_92792; // @[AxiLoadQueue.scala 246:86:@38344.8]
  wire  _T_92793; // @[AxiLoadQueue.scala 246:86:@38345.8]
  wire  _T_92794; // @[AxiLoadQueue.scala 246:86:@38346.8]
  wire  _T_92795; // @[AxiLoadQueue.scala 246:86:@38347.8]
  wire  _T_92796; // @[AxiLoadQueue.scala 246:86:@38348.8]
  wire  _T_92798; // @[AxiLoadQueue.scala 246:38:@38349.8]
  wire  _T_92817; // @[AxiLoadQueue.scala 247:11:@38366.8]
  wire  _T_92818; // @[AxiLoadQueue.scala 246:103:@38367.8]
  wire  _GEN_2020; // @[AxiLoadQueue.scala 243:104:@38332.6]
  wire  loadRequest_5; // @[AxiLoadQueue.scala 242:71:@38326.4]
  wire [15:0] _T_90472; // @[Mux.scala 31:69:@36525.4]
  wire  _T_92686; // @[AxiLoadQueue.scala 242:41:@38242.4]
  wire  _T_92687; // @[AxiLoadQueue.scala 242:38:@38243.4]
  wire  _T_92689; // @[AxiLoadQueue.scala 243:12:@38245.6]
  reg  loadInitiated_4; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_750;
  wire  _T_92691; // @[AxiLoadQueue.scala 243:46:@38246.6]
  wire  _T_92692; // @[AxiLoadQueue.scala 243:43:@38247.6]
  wire  _T_92694; // @[AxiLoadQueue.scala 243:78:@38248.6]
  wire  _T_92695; // @[AxiLoadQueue.scala 243:75:@38249.6]
  wire  _T_92698; // @[AxiLoadQueue.scala 246:86:@38252.8]
  wire  _T_92699; // @[AxiLoadQueue.scala 246:86:@38253.8]
  wire  _T_92700; // @[AxiLoadQueue.scala 246:86:@38254.8]
  wire  _T_92701; // @[AxiLoadQueue.scala 246:86:@38255.8]
  wire  _T_92702; // @[AxiLoadQueue.scala 246:86:@38256.8]
  wire  _T_92703; // @[AxiLoadQueue.scala 246:86:@38257.8]
  wire  _T_92704; // @[AxiLoadQueue.scala 246:86:@38258.8]
  wire  _T_92705; // @[AxiLoadQueue.scala 246:86:@38259.8]
  wire  _T_92706; // @[AxiLoadQueue.scala 246:86:@38260.8]
  wire  _T_92707; // @[AxiLoadQueue.scala 246:86:@38261.8]
  wire  _T_92708; // @[AxiLoadQueue.scala 246:86:@38262.8]
  wire  _T_92709; // @[AxiLoadQueue.scala 246:86:@38263.8]
  wire  _T_92710; // @[AxiLoadQueue.scala 246:86:@38264.8]
  wire  _T_92711; // @[AxiLoadQueue.scala 246:86:@38265.8]
  wire  _T_92712; // @[AxiLoadQueue.scala 246:86:@38266.8]
  wire  _T_92714; // @[AxiLoadQueue.scala 246:38:@38267.8]
  wire  _T_92733; // @[AxiLoadQueue.scala 247:11:@38284.8]
  wire  _T_92734; // @[AxiLoadQueue.scala 246:103:@38285.8]
  wire  _GEN_2016; // @[AxiLoadQueue.scala 243:104:@38250.6]
  wire  loadRequest_4; // @[AxiLoadQueue.scala 242:71:@38244.4]
  wire [15:0] _T_90473; // @[Mux.scala 31:69:@36526.4]
  wire  _T_92602; // @[AxiLoadQueue.scala 242:41:@38160.4]
  wire  _T_92603; // @[AxiLoadQueue.scala 242:38:@38161.4]
  wire  _T_92605; // @[AxiLoadQueue.scala 243:12:@38163.6]
  reg  loadInitiated_3; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_751;
  wire  _T_92607; // @[AxiLoadQueue.scala 243:46:@38164.6]
  wire  _T_92608; // @[AxiLoadQueue.scala 243:43:@38165.6]
  wire  _T_92610; // @[AxiLoadQueue.scala 243:78:@38166.6]
  wire  _T_92611; // @[AxiLoadQueue.scala 243:75:@38167.6]
  wire  _T_92614; // @[AxiLoadQueue.scala 246:86:@38170.8]
  wire  _T_92615; // @[AxiLoadQueue.scala 246:86:@38171.8]
  wire  _T_92616; // @[AxiLoadQueue.scala 246:86:@38172.8]
  wire  _T_92617; // @[AxiLoadQueue.scala 246:86:@38173.8]
  wire  _T_92618; // @[AxiLoadQueue.scala 246:86:@38174.8]
  wire  _T_92619; // @[AxiLoadQueue.scala 246:86:@38175.8]
  wire  _T_92620; // @[AxiLoadQueue.scala 246:86:@38176.8]
  wire  _T_92621; // @[AxiLoadQueue.scala 246:86:@38177.8]
  wire  _T_92622; // @[AxiLoadQueue.scala 246:86:@38178.8]
  wire  _T_92623; // @[AxiLoadQueue.scala 246:86:@38179.8]
  wire  _T_92624; // @[AxiLoadQueue.scala 246:86:@38180.8]
  wire  _T_92625; // @[AxiLoadQueue.scala 246:86:@38181.8]
  wire  _T_92626; // @[AxiLoadQueue.scala 246:86:@38182.8]
  wire  _T_92627; // @[AxiLoadQueue.scala 246:86:@38183.8]
  wire  _T_92628; // @[AxiLoadQueue.scala 246:86:@38184.8]
  wire  _T_92630; // @[AxiLoadQueue.scala 246:38:@38185.8]
  wire  _T_92649; // @[AxiLoadQueue.scala 247:11:@38202.8]
  wire  _T_92650; // @[AxiLoadQueue.scala 246:103:@38203.8]
  wire  _GEN_2012; // @[AxiLoadQueue.scala 243:104:@38168.6]
  wire  loadRequest_3; // @[AxiLoadQueue.scala 242:71:@38162.4]
  wire [15:0] _T_90474; // @[Mux.scala 31:69:@36527.4]
  wire  _T_92518; // @[AxiLoadQueue.scala 242:41:@38078.4]
  wire  _T_92519; // @[AxiLoadQueue.scala 242:38:@38079.4]
  wire  _T_92521; // @[AxiLoadQueue.scala 243:12:@38081.6]
  reg  loadInitiated_2; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_752;
  wire  _T_92523; // @[AxiLoadQueue.scala 243:46:@38082.6]
  wire  _T_92524; // @[AxiLoadQueue.scala 243:43:@38083.6]
  wire  _T_92526; // @[AxiLoadQueue.scala 243:78:@38084.6]
  wire  _T_92527; // @[AxiLoadQueue.scala 243:75:@38085.6]
  wire  _T_92530; // @[AxiLoadQueue.scala 246:86:@38088.8]
  wire  _T_92531; // @[AxiLoadQueue.scala 246:86:@38089.8]
  wire  _T_92532; // @[AxiLoadQueue.scala 246:86:@38090.8]
  wire  _T_92533; // @[AxiLoadQueue.scala 246:86:@38091.8]
  wire  _T_92534; // @[AxiLoadQueue.scala 246:86:@38092.8]
  wire  _T_92535; // @[AxiLoadQueue.scala 246:86:@38093.8]
  wire  _T_92536; // @[AxiLoadQueue.scala 246:86:@38094.8]
  wire  _T_92537; // @[AxiLoadQueue.scala 246:86:@38095.8]
  wire  _T_92538; // @[AxiLoadQueue.scala 246:86:@38096.8]
  wire  _T_92539; // @[AxiLoadQueue.scala 246:86:@38097.8]
  wire  _T_92540; // @[AxiLoadQueue.scala 246:86:@38098.8]
  wire  _T_92541; // @[AxiLoadQueue.scala 246:86:@38099.8]
  wire  _T_92542; // @[AxiLoadQueue.scala 246:86:@38100.8]
  wire  _T_92543; // @[AxiLoadQueue.scala 246:86:@38101.8]
  wire  _T_92544; // @[AxiLoadQueue.scala 246:86:@38102.8]
  wire  _T_92546; // @[AxiLoadQueue.scala 246:38:@38103.8]
  wire  _T_92565; // @[AxiLoadQueue.scala 247:11:@38120.8]
  wire  _T_92566; // @[AxiLoadQueue.scala 246:103:@38121.8]
  wire  _GEN_2008; // @[AxiLoadQueue.scala 243:104:@38086.6]
  wire  loadRequest_2; // @[AxiLoadQueue.scala 242:71:@38080.4]
  wire [15:0] _T_90475; // @[Mux.scala 31:69:@36528.4]
  wire  _T_92434; // @[AxiLoadQueue.scala 242:41:@37996.4]
  wire  _T_92435; // @[AxiLoadQueue.scala 242:38:@37997.4]
  wire  _T_92437; // @[AxiLoadQueue.scala 243:12:@37999.6]
  reg  loadInitiated_1; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_753;
  wire  _T_92439; // @[AxiLoadQueue.scala 243:46:@38000.6]
  wire  _T_92440; // @[AxiLoadQueue.scala 243:43:@38001.6]
  wire  _T_92442; // @[AxiLoadQueue.scala 243:78:@38002.6]
  wire  _T_92443; // @[AxiLoadQueue.scala 243:75:@38003.6]
  wire  _T_92446; // @[AxiLoadQueue.scala 246:86:@38006.8]
  wire  _T_92447; // @[AxiLoadQueue.scala 246:86:@38007.8]
  wire  _T_92448; // @[AxiLoadQueue.scala 246:86:@38008.8]
  wire  _T_92449; // @[AxiLoadQueue.scala 246:86:@38009.8]
  wire  _T_92450; // @[AxiLoadQueue.scala 246:86:@38010.8]
  wire  _T_92451; // @[AxiLoadQueue.scala 246:86:@38011.8]
  wire  _T_92452; // @[AxiLoadQueue.scala 246:86:@38012.8]
  wire  _T_92453; // @[AxiLoadQueue.scala 246:86:@38013.8]
  wire  _T_92454; // @[AxiLoadQueue.scala 246:86:@38014.8]
  wire  _T_92455; // @[AxiLoadQueue.scala 246:86:@38015.8]
  wire  _T_92456; // @[AxiLoadQueue.scala 246:86:@38016.8]
  wire  _T_92457; // @[AxiLoadQueue.scala 246:86:@38017.8]
  wire  _T_92458; // @[AxiLoadQueue.scala 246:86:@38018.8]
  wire  _T_92459; // @[AxiLoadQueue.scala 246:86:@38019.8]
  wire  _T_92460; // @[AxiLoadQueue.scala 246:86:@38020.8]
  wire  _T_92462; // @[AxiLoadQueue.scala 246:38:@38021.8]
  wire  _T_92481; // @[AxiLoadQueue.scala 247:11:@38038.8]
  wire  _T_92482; // @[AxiLoadQueue.scala 246:103:@38039.8]
  wire  _GEN_2004; // @[AxiLoadQueue.scala 243:104:@38004.6]
  wire  loadRequest_1; // @[AxiLoadQueue.scala 242:71:@37998.4]
  wire [15:0] _T_90476; // @[Mux.scala 31:69:@36529.4]
  wire  _T_92350; // @[AxiLoadQueue.scala 242:41:@37914.4]
  wire  _T_92351; // @[AxiLoadQueue.scala 242:38:@37915.4]
  wire  _T_92353; // @[AxiLoadQueue.scala 243:12:@37917.6]
  reg  loadInitiated_0; // @[AxiLoadQueue.scala 207:30:@37622.4]
  reg [31:0] _RAND_754;
  wire  _T_92355; // @[AxiLoadQueue.scala 243:46:@37918.6]
  wire  _T_92356; // @[AxiLoadQueue.scala 243:43:@37919.6]
  wire  _T_92358; // @[AxiLoadQueue.scala 243:78:@37920.6]
  wire  _T_92359; // @[AxiLoadQueue.scala 243:75:@37921.6]
  wire  _T_92362; // @[AxiLoadQueue.scala 246:86:@37924.8]
  wire  _T_92363; // @[AxiLoadQueue.scala 246:86:@37925.8]
  wire  _T_92364; // @[AxiLoadQueue.scala 246:86:@37926.8]
  wire  _T_92365; // @[AxiLoadQueue.scala 246:86:@37927.8]
  wire  _T_92366; // @[AxiLoadQueue.scala 246:86:@37928.8]
  wire  _T_92367; // @[AxiLoadQueue.scala 246:86:@37929.8]
  wire  _T_92368; // @[AxiLoadQueue.scala 246:86:@37930.8]
  wire  _T_92369; // @[AxiLoadQueue.scala 246:86:@37931.8]
  wire  _T_92370; // @[AxiLoadQueue.scala 246:86:@37932.8]
  wire  _T_92371; // @[AxiLoadQueue.scala 246:86:@37933.8]
  wire  _T_92372; // @[AxiLoadQueue.scala 246:86:@37934.8]
  wire  _T_92373; // @[AxiLoadQueue.scala 246:86:@37935.8]
  wire  _T_92374; // @[AxiLoadQueue.scala 246:86:@37936.8]
  wire  _T_92375; // @[AxiLoadQueue.scala 246:86:@37937.8]
  wire  _T_92376; // @[AxiLoadQueue.scala 246:86:@37938.8]
  wire  _T_92378; // @[AxiLoadQueue.scala 246:38:@37939.8]
  wire  _T_92397; // @[AxiLoadQueue.scala 247:11:@37956.8]
  wire  _T_92398; // @[AxiLoadQueue.scala 246:103:@37957.8]
  wire  _GEN_2000; // @[AxiLoadQueue.scala 243:104:@37922.6]
  wire  loadRequest_0; // @[AxiLoadQueue.scala 242:71:@37916.4]
  wire [15:0] _T_90477; // @[Mux.scala 31:69:@36530.4]
  wire  _T_90478; // @[OneHot.scala 66:30:@36531.4]
  wire  _T_90479; // @[OneHot.scala 66:30:@36532.4]
  wire  _T_90480; // @[OneHot.scala 66:30:@36533.4]
  wire  _T_90481; // @[OneHot.scala 66:30:@36534.4]
  wire  _T_90482; // @[OneHot.scala 66:30:@36535.4]
  wire  _T_90483; // @[OneHot.scala 66:30:@36536.4]
  wire  _T_90484; // @[OneHot.scala 66:30:@36537.4]
  wire  _T_90485; // @[OneHot.scala 66:30:@36538.4]
  wire  _T_90486; // @[OneHot.scala 66:30:@36539.4]
  wire  _T_90487; // @[OneHot.scala 66:30:@36540.4]
  wire  _T_90488; // @[OneHot.scala 66:30:@36541.4]
  wire  _T_90489; // @[OneHot.scala 66:30:@36542.4]
  wire  _T_90490; // @[OneHot.scala 66:30:@36543.4]
  wire  _T_90491; // @[OneHot.scala 66:30:@36544.4]
  wire  _T_90492; // @[OneHot.scala 66:30:@36545.4]
  wire  _T_90493; // @[OneHot.scala 66:30:@36546.4]
  wire [15:0] _T_90534; // @[Mux.scala 31:69:@36564.4]
  wire [15:0] _T_90535; // @[Mux.scala 31:69:@36565.4]
  wire [15:0] _T_90536; // @[Mux.scala 31:69:@36566.4]
  wire [15:0] _T_90537; // @[Mux.scala 31:69:@36567.4]
  wire [15:0] _T_90538; // @[Mux.scala 31:69:@36568.4]
  wire [15:0] _T_90539; // @[Mux.scala 31:69:@36569.4]
  wire [15:0] _T_90540; // @[Mux.scala 31:69:@36570.4]
  wire [15:0] _T_90541; // @[Mux.scala 31:69:@36571.4]
  wire [15:0] _T_90542; // @[Mux.scala 31:69:@36572.4]
  wire [15:0] _T_90543; // @[Mux.scala 31:69:@36573.4]
  wire [15:0] _T_90544; // @[Mux.scala 31:69:@36574.4]
  wire [15:0] _T_90545; // @[Mux.scala 31:69:@36575.4]
  wire [15:0] _T_90546; // @[Mux.scala 31:69:@36576.4]
  wire [15:0] _T_90547; // @[Mux.scala 31:69:@36577.4]
  wire [15:0] _T_90548; // @[Mux.scala 31:69:@36578.4]
  wire [15:0] _T_90549; // @[Mux.scala 31:69:@36579.4]
  wire  _T_90550; // @[OneHot.scala 66:30:@36580.4]
  wire  _T_90551; // @[OneHot.scala 66:30:@36581.4]
  wire  _T_90552; // @[OneHot.scala 66:30:@36582.4]
  wire  _T_90553; // @[OneHot.scala 66:30:@36583.4]
  wire  _T_90554; // @[OneHot.scala 66:30:@36584.4]
  wire  _T_90555; // @[OneHot.scala 66:30:@36585.4]
  wire  _T_90556; // @[OneHot.scala 66:30:@36586.4]
  wire  _T_90557; // @[OneHot.scala 66:30:@36587.4]
  wire  _T_90558; // @[OneHot.scala 66:30:@36588.4]
  wire  _T_90559; // @[OneHot.scala 66:30:@36589.4]
  wire  _T_90560; // @[OneHot.scala 66:30:@36590.4]
  wire  _T_90561; // @[OneHot.scala 66:30:@36591.4]
  wire  _T_90562; // @[OneHot.scala 66:30:@36592.4]
  wire  _T_90563; // @[OneHot.scala 66:30:@36593.4]
  wire  _T_90564; // @[OneHot.scala 66:30:@36594.4]
  wire  _T_90565; // @[OneHot.scala 66:30:@36595.4]
  wire [15:0] _T_90606; // @[Mux.scala 31:69:@36613.4]
  wire [15:0] _T_90607; // @[Mux.scala 31:69:@36614.4]
  wire [15:0] _T_90608; // @[Mux.scala 31:69:@36615.4]
  wire [15:0] _T_90609; // @[Mux.scala 31:69:@36616.4]
  wire [15:0] _T_90610; // @[Mux.scala 31:69:@36617.4]
  wire [15:0] _T_90611; // @[Mux.scala 31:69:@36618.4]
  wire [15:0] _T_90612; // @[Mux.scala 31:69:@36619.4]
  wire [15:0] _T_90613; // @[Mux.scala 31:69:@36620.4]
  wire [15:0] _T_90614; // @[Mux.scala 31:69:@36621.4]
  wire [15:0] _T_90615; // @[Mux.scala 31:69:@36622.4]
  wire [15:0] _T_90616; // @[Mux.scala 31:69:@36623.4]
  wire [15:0] _T_90617; // @[Mux.scala 31:69:@36624.4]
  wire [15:0] _T_90618; // @[Mux.scala 31:69:@36625.4]
  wire [15:0] _T_90619; // @[Mux.scala 31:69:@36626.4]
  wire [15:0] _T_90620; // @[Mux.scala 31:69:@36627.4]
  wire [15:0] _T_90621; // @[Mux.scala 31:69:@36628.4]
  wire  _T_90622; // @[OneHot.scala 66:30:@36629.4]
  wire  _T_90623; // @[OneHot.scala 66:30:@36630.4]
  wire  _T_90624; // @[OneHot.scala 66:30:@36631.4]
  wire  _T_90625; // @[OneHot.scala 66:30:@36632.4]
  wire  _T_90626; // @[OneHot.scala 66:30:@36633.4]
  wire  _T_90627; // @[OneHot.scala 66:30:@36634.4]
  wire  _T_90628; // @[OneHot.scala 66:30:@36635.4]
  wire  _T_90629; // @[OneHot.scala 66:30:@36636.4]
  wire  _T_90630; // @[OneHot.scala 66:30:@36637.4]
  wire  _T_90631; // @[OneHot.scala 66:30:@36638.4]
  wire  _T_90632; // @[OneHot.scala 66:30:@36639.4]
  wire  _T_90633; // @[OneHot.scala 66:30:@36640.4]
  wire  _T_90634; // @[OneHot.scala 66:30:@36641.4]
  wire  _T_90635; // @[OneHot.scala 66:30:@36642.4]
  wire  _T_90636; // @[OneHot.scala 66:30:@36643.4]
  wire  _T_90637; // @[OneHot.scala 66:30:@36644.4]
  wire [15:0] _T_90678; // @[Mux.scala 31:69:@36662.4]
  wire [15:0] _T_90679; // @[Mux.scala 31:69:@36663.4]
  wire [15:0] _T_90680; // @[Mux.scala 31:69:@36664.4]
  wire [15:0] _T_90681; // @[Mux.scala 31:69:@36665.4]
  wire [15:0] _T_90682; // @[Mux.scala 31:69:@36666.4]
  wire [15:0] _T_90683; // @[Mux.scala 31:69:@36667.4]
  wire [15:0] _T_90684; // @[Mux.scala 31:69:@36668.4]
  wire [15:0] _T_90685; // @[Mux.scala 31:69:@36669.4]
  wire [15:0] _T_90686; // @[Mux.scala 31:69:@36670.4]
  wire [15:0] _T_90687; // @[Mux.scala 31:69:@36671.4]
  wire [15:0] _T_90688; // @[Mux.scala 31:69:@36672.4]
  wire [15:0] _T_90689; // @[Mux.scala 31:69:@36673.4]
  wire [15:0] _T_90690; // @[Mux.scala 31:69:@36674.4]
  wire [15:0] _T_90691; // @[Mux.scala 31:69:@36675.4]
  wire [15:0] _T_90692; // @[Mux.scala 31:69:@36676.4]
  wire [15:0] _T_90693; // @[Mux.scala 31:69:@36677.4]
  wire  _T_90694; // @[OneHot.scala 66:30:@36678.4]
  wire  _T_90695; // @[OneHot.scala 66:30:@36679.4]
  wire  _T_90696; // @[OneHot.scala 66:30:@36680.4]
  wire  _T_90697; // @[OneHot.scala 66:30:@36681.4]
  wire  _T_90698; // @[OneHot.scala 66:30:@36682.4]
  wire  _T_90699; // @[OneHot.scala 66:30:@36683.4]
  wire  _T_90700; // @[OneHot.scala 66:30:@36684.4]
  wire  _T_90701; // @[OneHot.scala 66:30:@36685.4]
  wire  _T_90702; // @[OneHot.scala 66:30:@36686.4]
  wire  _T_90703; // @[OneHot.scala 66:30:@36687.4]
  wire  _T_90704; // @[OneHot.scala 66:30:@36688.4]
  wire  _T_90705; // @[OneHot.scala 66:30:@36689.4]
  wire  _T_90706; // @[OneHot.scala 66:30:@36690.4]
  wire  _T_90707; // @[OneHot.scala 66:30:@36691.4]
  wire  _T_90708; // @[OneHot.scala 66:30:@36692.4]
  wire  _T_90709; // @[OneHot.scala 66:30:@36693.4]
  wire [15:0] _T_90750; // @[Mux.scala 31:69:@36711.4]
  wire [15:0] _T_90751; // @[Mux.scala 31:69:@36712.4]
  wire [15:0] _T_90752; // @[Mux.scala 31:69:@36713.4]
  wire [15:0] _T_90753; // @[Mux.scala 31:69:@36714.4]
  wire [15:0] _T_90754; // @[Mux.scala 31:69:@36715.4]
  wire [15:0] _T_90755; // @[Mux.scala 31:69:@36716.4]
  wire [15:0] _T_90756; // @[Mux.scala 31:69:@36717.4]
  wire [15:0] _T_90757; // @[Mux.scala 31:69:@36718.4]
  wire [15:0] _T_90758; // @[Mux.scala 31:69:@36719.4]
  wire [15:0] _T_90759; // @[Mux.scala 31:69:@36720.4]
  wire [15:0] _T_90760; // @[Mux.scala 31:69:@36721.4]
  wire [15:0] _T_90761; // @[Mux.scala 31:69:@36722.4]
  wire [15:0] _T_90762; // @[Mux.scala 31:69:@36723.4]
  wire [15:0] _T_90763; // @[Mux.scala 31:69:@36724.4]
  wire [15:0] _T_90764; // @[Mux.scala 31:69:@36725.4]
  wire [15:0] _T_90765; // @[Mux.scala 31:69:@36726.4]
  wire  _T_90766; // @[OneHot.scala 66:30:@36727.4]
  wire  _T_90767; // @[OneHot.scala 66:30:@36728.4]
  wire  _T_90768; // @[OneHot.scala 66:30:@36729.4]
  wire  _T_90769; // @[OneHot.scala 66:30:@36730.4]
  wire  _T_90770; // @[OneHot.scala 66:30:@36731.4]
  wire  _T_90771; // @[OneHot.scala 66:30:@36732.4]
  wire  _T_90772; // @[OneHot.scala 66:30:@36733.4]
  wire  _T_90773; // @[OneHot.scala 66:30:@36734.4]
  wire  _T_90774; // @[OneHot.scala 66:30:@36735.4]
  wire  _T_90775; // @[OneHot.scala 66:30:@36736.4]
  wire  _T_90776; // @[OneHot.scala 66:30:@36737.4]
  wire  _T_90777; // @[OneHot.scala 66:30:@36738.4]
  wire  _T_90778; // @[OneHot.scala 66:30:@36739.4]
  wire  _T_90779; // @[OneHot.scala 66:30:@36740.4]
  wire  _T_90780; // @[OneHot.scala 66:30:@36741.4]
  wire  _T_90781; // @[OneHot.scala 66:30:@36742.4]
  wire [15:0] _T_90822; // @[Mux.scala 31:69:@36760.4]
  wire [15:0] _T_90823; // @[Mux.scala 31:69:@36761.4]
  wire [15:0] _T_90824; // @[Mux.scala 31:69:@36762.4]
  wire [15:0] _T_90825; // @[Mux.scala 31:69:@36763.4]
  wire [15:0] _T_90826; // @[Mux.scala 31:69:@36764.4]
  wire [15:0] _T_90827; // @[Mux.scala 31:69:@36765.4]
  wire [15:0] _T_90828; // @[Mux.scala 31:69:@36766.4]
  wire [15:0] _T_90829; // @[Mux.scala 31:69:@36767.4]
  wire [15:0] _T_90830; // @[Mux.scala 31:69:@36768.4]
  wire [15:0] _T_90831; // @[Mux.scala 31:69:@36769.4]
  wire [15:0] _T_90832; // @[Mux.scala 31:69:@36770.4]
  wire [15:0] _T_90833; // @[Mux.scala 31:69:@36771.4]
  wire [15:0] _T_90834; // @[Mux.scala 31:69:@36772.4]
  wire [15:0] _T_90835; // @[Mux.scala 31:69:@36773.4]
  wire [15:0] _T_90836; // @[Mux.scala 31:69:@36774.4]
  wire [15:0] _T_90837; // @[Mux.scala 31:69:@36775.4]
  wire  _T_90838; // @[OneHot.scala 66:30:@36776.4]
  wire  _T_90839; // @[OneHot.scala 66:30:@36777.4]
  wire  _T_90840; // @[OneHot.scala 66:30:@36778.4]
  wire  _T_90841; // @[OneHot.scala 66:30:@36779.4]
  wire  _T_90842; // @[OneHot.scala 66:30:@36780.4]
  wire  _T_90843; // @[OneHot.scala 66:30:@36781.4]
  wire  _T_90844; // @[OneHot.scala 66:30:@36782.4]
  wire  _T_90845; // @[OneHot.scala 66:30:@36783.4]
  wire  _T_90846; // @[OneHot.scala 66:30:@36784.4]
  wire  _T_90847; // @[OneHot.scala 66:30:@36785.4]
  wire  _T_90848; // @[OneHot.scala 66:30:@36786.4]
  wire  _T_90849; // @[OneHot.scala 66:30:@36787.4]
  wire  _T_90850; // @[OneHot.scala 66:30:@36788.4]
  wire  _T_90851; // @[OneHot.scala 66:30:@36789.4]
  wire  _T_90852; // @[OneHot.scala 66:30:@36790.4]
  wire  _T_90853; // @[OneHot.scala 66:30:@36791.4]
  wire [15:0] _T_90894; // @[Mux.scala 31:69:@36809.4]
  wire [15:0] _T_90895; // @[Mux.scala 31:69:@36810.4]
  wire [15:0] _T_90896; // @[Mux.scala 31:69:@36811.4]
  wire [15:0] _T_90897; // @[Mux.scala 31:69:@36812.4]
  wire [15:0] _T_90898; // @[Mux.scala 31:69:@36813.4]
  wire [15:0] _T_90899; // @[Mux.scala 31:69:@36814.4]
  wire [15:0] _T_90900; // @[Mux.scala 31:69:@36815.4]
  wire [15:0] _T_90901; // @[Mux.scala 31:69:@36816.4]
  wire [15:0] _T_90902; // @[Mux.scala 31:69:@36817.4]
  wire [15:0] _T_90903; // @[Mux.scala 31:69:@36818.4]
  wire [15:0] _T_90904; // @[Mux.scala 31:69:@36819.4]
  wire [15:0] _T_90905; // @[Mux.scala 31:69:@36820.4]
  wire [15:0] _T_90906; // @[Mux.scala 31:69:@36821.4]
  wire [15:0] _T_90907; // @[Mux.scala 31:69:@36822.4]
  wire [15:0] _T_90908; // @[Mux.scala 31:69:@36823.4]
  wire [15:0] _T_90909; // @[Mux.scala 31:69:@36824.4]
  wire  _T_90910; // @[OneHot.scala 66:30:@36825.4]
  wire  _T_90911; // @[OneHot.scala 66:30:@36826.4]
  wire  _T_90912; // @[OneHot.scala 66:30:@36827.4]
  wire  _T_90913; // @[OneHot.scala 66:30:@36828.4]
  wire  _T_90914; // @[OneHot.scala 66:30:@36829.4]
  wire  _T_90915; // @[OneHot.scala 66:30:@36830.4]
  wire  _T_90916; // @[OneHot.scala 66:30:@36831.4]
  wire  _T_90917; // @[OneHot.scala 66:30:@36832.4]
  wire  _T_90918; // @[OneHot.scala 66:30:@36833.4]
  wire  _T_90919; // @[OneHot.scala 66:30:@36834.4]
  wire  _T_90920; // @[OneHot.scala 66:30:@36835.4]
  wire  _T_90921; // @[OneHot.scala 66:30:@36836.4]
  wire  _T_90922; // @[OneHot.scala 66:30:@36837.4]
  wire  _T_90923; // @[OneHot.scala 66:30:@36838.4]
  wire  _T_90924; // @[OneHot.scala 66:30:@36839.4]
  wire  _T_90925; // @[OneHot.scala 66:30:@36840.4]
  wire [15:0] _T_90966; // @[Mux.scala 31:69:@36858.4]
  wire [15:0] _T_90967; // @[Mux.scala 31:69:@36859.4]
  wire [15:0] _T_90968; // @[Mux.scala 31:69:@36860.4]
  wire [15:0] _T_90969; // @[Mux.scala 31:69:@36861.4]
  wire [15:0] _T_90970; // @[Mux.scala 31:69:@36862.4]
  wire [15:0] _T_90971; // @[Mux.scala 31:69:@36863.4]
  wire [15:0] _T_90972; // @[Mux.scala 31:69:@36864.4]
  wire [15:0] _T_90973; // @[Mux.scala 31:69:@36865.4]
  wire [15:0] _T_90974; // @[Mux.scala 31:69:@36866.4]
  wire [15:0] _T_90975; // @[Mux.scala 31:69:@36867.4]
  wire [15:0] _T_90976; // @[Mux.scala 31:69:@36868.4]
  wire [15:0] _T_90977; // @[Mux.scala 31:69:@36869.4]
  wire [15:0] _T_90978; // @[Mux.scala 31:69:@36870.4]
  wire [15:0] _T_90979; // @[Mux.scala 31:69:@36871.4]
  wire [15:0] _T_90980; // @[Mux.scala 31:69:@36872.4]
  wire [15:0] _T_90981; // @[Mux.scala 31:69:@36873.4]
  wire  _T_90982; // @[OneHot.scala 66:30:@36874.4]
  wire  _T_90983; // @[OneHot.scala 66:30:@36875.4]
  wire  _T_90984; // @[OneHot.scala 66:30:@36876.4]
  wire  _T_90985; // @[OneHot.scala 66:30:@36877.4]
  wire  _T_90986; // @[OneHot.scala 66:30:@36878.4]
  wire  _T_90987; // @[OneHot.scala 66:30:@36879.4]
  wire  _T_90988; // @[OneHot.scala 66:30:@36880.4]
  wire  _T_90989; // @[OneHot.scala 66:30:@36881.4]
  wire  _T_90990; // @[OneHot.scala 66:30:@36882.4]
  wire  _T_90991; // @[OneHot.scala 66:30:@36883.4]
  wire  _T_90992; // @[OneHot.scala 66:30:@36884.4]
  wire  _T_90993; // @[OneHot.scala 66:30:@36885.4]
  wire  _T_90994; // @[OneHot.scala 66:30:@36886.4]
  wire  _T_90995; // @[OneHot.scala 66:30:@36887.4]
  wire  _T_90996; // @[OneHot.scala 66:30:@36888.4]
  wire  _T_90997; // @[OneHot.scala 66:30:@36889.4]
  wire [15:0] _T_91038; // @[Mux.scala 31:69:@36907.4]
  wire [15:0] _T_91039; // @[Mux.scala 31:69:@36908.4]
  wire [15:0] _T_91040; // @[Mux.scala 31:69:@36909.4]
  wire [15:0] _T_91041; // @[Mux.scala 31:69:@36910.4]
  wire [15:0] _T_91042; // @[Mux.scala 31:69:@36911.4]
  wire [15:0] _T_91043; // @[Mux.scala 31:69:@36912.4]
  wire [15:0] _T_91044; // @[Mux.scala 31:69:@36913.4]
  wire [15:0] _T_91045; // @[Mux.scala 31:69:@36914.4]
  wire [15:0] _T_91046; // @[Mux.scala 31:69:@36915.4]
  wire [15:0] _T_91047; // @[Mux.scala 31:69:@36916.4]
  wire [15:0] _T_91048; // @[Mux.scala 31:69:@36917.4]
  wire [15:0] _T_91049; // @[Mux.scala 31:69:@36918.4]
  wire [15:0] _T_91050; // @[Mux.scala 31:69:@36919.4]
  wire [15:0] _T_91051; // @[Mux.scala 31:69:@36920.4]
  wire [15:0] _T_91052; // @[Mux.scala 31:69:@36921.4]
  wire [15:0] _T_91053; // @[Mux.scala 31:69:@36922.4]
  wire  _T_91054; // @[OneHot.scala 66:30:@36923.4]
  wire  _T_91055; // @[OneHot.scala 66:30:@36924.4]
  wire  _T_91056; // @[OneHot.scala 66:30:@36925.4]
  wire  _T_91057; // @[OneHot.scala 66:30:@36926.4]
  wire  _T_91058; // @[OneHot.scala 66:30:@36927.4]
  wire  _T_91059; // @[OneHot.scala 66:30:@36928.4]
  wire  _T_91060; // @[OneHot.scala 66:30:@36929.4]
  wire  _T_91061; // @[OneHot.scala 66:30:@36930.4]
  wire  _T_91062; // @[OneHot.scala 66:30:@36931.4]
  wire  _T_91063; // @[OneHot.scala 66:30:@36932.4]
  wire  _T_91064; // @[OneHot.scala 66:30:@36933.4]
  wire  _T_91065; // @[OneHot.scala 66:30:@36934.4]
  wire  _T_91066; // @[OneHot.scala 66:30:@36935.4]
  wire  _T_91067; // @[OneHot.scala 66:30:@36936.4]
  wire  _T_91068; // @[OneHot.scala 66:30:@36937.4]
  wire  _T_91069; // @[OneHot.scala 66:30:@36938.4]
  wire [15:0] _T_91110; // @[Mux.scala 31:69:@36956.4]
  wire [15:0] _T_91111; // @[Mux.scala 31:69:@36957.4]
  wire [15:0] _T_91112; // @[Mux.scala 31:69:@36958.4]
  wire [15:0] _T_91113; // @[Mux.scala 31:69:@36959.4]
  wire [15:0] _T_91114; // @[Mux.scala 31:69:@36960.4]
  wire [15:0] _T_91115; // @[Mux.scala 31:69:@36961.4]
  wire [15:0] _T_91116; // @[Mux.scala 31:69:@36962.4]
  wire [15:0] _T_91117; // @[Mux.scala 31:69:@36963.4]
  wire [15:0] _T_91118; // @[Mux.scala 31:69:@36964.4]
  wire [15:0] _T_91119; // @[Mux.scala 31:69:@36965.4]
  wire [15:0] _T_91120; // @[Mux.scala 31:69:@36966.4]
  wire [15:0] _T_91121; // @[Mux.scala 31:69:@36967.4]
  wire [15:0] _T_91122; // @[Mux.scala 31:69:@36968.4]
  wire [15:0] _T_91123; // @[Mux.scala 31:69:@36969.4]
  wire [15:0] _T_91124; // @[Mux.scala 31:69:@36970.4]
  wire [15:0] _T_91125; // @[Mux.scala 31:69:@36971.4]
  wire  _T_91126; // @[OneHot.scala 66:30:@36972.4]
  wire  _T_91127; // @[OneHot.scala 66:30:@36973.4]
  wire  _T_91128; // @[OneHot.scala 66:30:@36974.4]
  wire  _T_91129; // @[OneHot.scala 66:30:@36975.4]
  wire  _T_91130; // @[OneHot.scala 66:30:@36976.4]
  wire  _T_91131; // @[OneHot.scala 66:30:@36977.4]
  wire  _T_91132; // @[OneHot.scala 66:30:@36978.4]
  wire  _T_91133; // @[OneHot.scala 66:30:@36979.4]
  wire  _T_91134; // @[OneHot.scala 66:30:@36980.4]
  wire  _T_91135; // @[OneHot.scala 66:30:@36981.4]
  wire  _T_91136; // @[OneHot.scala 66:30:@36982.4]
  wire  _T_91137; // @[OneHot.scala 66:30:@36983.4]
  wire  _T_91138; // @[OneHot.scala 66:30:@36984.4]
  wire  _T_91139; // @[OneHot.scala 66:30:@36985.4]
  wire  _T_91140; // @[OneHot.scala 66:30:@36986.4]
  wire  _T_91141; // @[OneHot.scala 66:30:@36987.4]
  wire [15:0] _T_91182; // @[Mux.scala 31:69:@37005.4]
  wire [15:0] _T_91183; // @[Mux.scala 31:69:@37006.4]
  wire [15:0] _T_91184; // @[Mux.scala 31:69:@37007.4]
  wire [15:0] _T_91185; // @[Mux.scala 31:69:@37008.4]
  wire [15:0] _T_91186; // @[Mux.scala 31:69:@37009.4]
  wire [15:0] _T_91187; // @[Mux.scala 31:69:@37010.4]
  wire [15:0] _T_91188; // @[Mux.scala 31:69:@37011.4]
  wire [15:0] _T_91189; // @[Mux.scala 31:69:@37012.4]
  wire [15:0] _T_91190; // @[Mux.scala 31:69:@37013.4]
  wire [15:0] _T_91191; // @[Mux.scala 31:69:@37014.4]
  wire [15:0] _T_91192; // @[Mux.scala 31:69:@37015.4]
  wire [15:0] _T_91193; // @[Mux.scala 31:69:@37016.4]
  wire [15:0] _T_91194; // @[Mux.scala 31:69:@37017.4]
  wire [15:0] _T_91195; // @[Mux.scala 31:69:@37018.4]
  wire [15:0] _T_91196; // @[Mux.scala 31:69:@37019.4]
  wire [15:0] _T_91197; // @[Mux.scala 31:69:@37020.4]
  wire  _T_91198; // @[OneHot.scala 66:30:@37021.4]
  wire  _T_91199; // @[OneHot.scala 66:30:@37022.4]
  wire  _T_91200; // @[OneHot.scala 66:30:@37023.4]
  wire  _T_91201; // @[OneHot.scala 66:30:@37024.4]
  wire  _T_91202; // @[OneHot.scala 66:30:@37025.4]
  wire  _T_91203; // @[OneHot.scala 66:30:@37026.4]
  wire  _T_91204; // @[OneHot.scala 66:30:@37027.4]
  wire  _T_91205; // @[OneHot.scala 66:30:@37028.4]
  wire  _T_91206; // @[OneHot.scala 66:30:@37029.4]
  wire  _T_91207; // @[OneHot.scala 66:30:@37030.4]
  wire  _T_91208; // @[OneHot.scala 66:30:@37031.4]
  wire  _T_91209; // @[OneHot.scala 66:30:@37032.4]
  wire  _T_91210; // @[OneHot.scala 66:30:@37033.4]
  wire  _T_91211; // @[OneHot.scala 66:30:@37034.4]
  wire  _T_91212; // @[OneHot.scala 66:30:@37035.4]
  wire  _T_91213; // @[OneHot.scala 66:30:@37036.4]
  wire [15:0] _T_91254; // @[Mux.scala 31:69:@37054.4]
  wire [15:0] _T_91255; // @[Mux.scala 31:69:@37055.4]
  wire [15:0] _T_91256; // @[Mux.scala 31:69:@37056.4]
  wire [15:0] _T_91257; // @[Mux.scala 31:69:@37057.4]
  wire [15:0] _T_91258; // @[Mux.scala 31:69:@37058.4]
  wire [15:0] _T_91259; // @[Mux.scala 31:69:@37059.4]
  wire [15:0] _T_91260; // @[Mux.scala 31:69:@37060.4]
  wire [15:0] _T_91261; // @[Mux.scala 31:69:@37061.4]
  wire [15:0] _T_91262; // @[Mux.scala 31:69:@37062.4]
  wire [15:0] _T_91263; // @[Mux.scala 31:69:@37063.4]
  wire [15:0] _T_91264; // @[Mux.scala 31:69:@37064.4]
  wire [15:0] _T_91265; // @[Mux.scala 31:69:@37065.4]
  wire [15:0] _T_91266; // @[Mux.scala 31:69:@37066.4]
  wire [15:0] _T_91267; // @[Mux.scala 31:69:@37067.4]
  wire [15:0] _T_91268; // @[Mux.scala 31:69:@37068.4]
  wire [15:0] _T_91269; // @[Mux.scala 31:69:@37069.4]
  wire  _T_91270; // @[OneHot.scala 66:30:@37070.4]
  wire  _T_91271; // @[OneHot.scala 66:30:@37071.4]
  wire  _T_91272; // @[OneHot.scala 66:30:@37072.4]
  wire  _T_91273; // @[OneHot.scala 66:30:@37073.4]
  wire  _T_91274; // @[OneHot.scala 66:30:@37074.4]
  wire  _T_91275; // @[OneHot.scala 66:30:@37075.4]
  wire  _T_91276; // @[OneHot.scala 66:30:@37076.4]
  wire  _T_91277; // @[OneHot.scala 66:30:@37077.4]
  wire  _T_91278; // @[OneHot.scala 66:30:@37078.4]
  wire  _T_91279; // @[OneHot.scala 66:30:@37079.4]
  wire  _T_91280; // @[OneHot.scala 66:30:@37080.4]
  wire  _T_91281; // @[OneHot.scala 66:30:@37081.4]
  wire  _T_91282; // @[OneHot.scala 66:30:@37082.4]
  wire  _T_91283; // @[OneHot.scala 66:30:@37083.4]
  wire  _T_91284; // @[OneHot.scala 66:30:@37084.4]
  wire  _T_91285; // @[OneHot.scala 66:30:@37085.4]
  wire [15:0] _T_91326; // @[Mux.scala 31:69:@37103.4]
  wire [15:0] _T_91327; // @[Mux.scala 31:69:@37104.4]
  wire [15:0] _T_91328; // @[Mux.scala 31:69:@37105.4]
  wire [15:0] _T_91329; // @[Mux.scala 31:69:@37106.4]
  wire [15:0] _T_91330; // @[Mux.scala 31:69:@37107.4]
  wire [15:0] _T_91331; // @[Mux.scala 31:69:@37108.4]
  wire [15:0] _T_91332; // @[Mux.scala 31:69:@37109.4]
  wire [15:0] _T_91333; // @[Mux.scala 31:69:@37110.4]
  wire [15:0] _T_91334; // @[Mux.scala 31:69:@37111.4]
  wire [15:0] _T_91335; // @[Mux.scala 31:69:@37112.4]
  wire [15:0] _T_91336; // @[Mux.scala 31:69:@37113.4]
  wire [15:0] _T_91337; // @[Mux.scala 31:69:@37114.4]
  wire [15:0] _T_91338; // @[Mux.scala 31:69:@37115.4]
  wire [15:0] _T_91339; // @[Mux.scala 31:69:@37116.4]
  wire [15:0] _T_91340; // @[Mux.scala 31:69:@37117.4]
  wire [15:0] _T_91341; // @[Mux.scala 31:69:@37118.4]
  wire  _T_91342; // @[OneHot.scala 66:30:@37119.4]
  wire  _T_91343; // @[OneHot.scala 66:30:@37120.4]
  wire  _T_91344; // @[OneHot.scala 66:30:@37121.4]
  wire  _T_91345; // @[OneHot.scala 66:30:@37122.4]
  wire  _T_91346; // @[OneHot.scala 66:30:@37123.4]
  wire  _T_91347; // @[OneHot.scala 66:30:@37124.4]
  wire  _T_91348; // @[OneHot.scala 66:30:@37125.4]
  wire  _T_91349; // @[OneHot.scala 66:30:@37126.4]
  wire  _T_91350; // @[OneHot.scala 66:30:@37127.4]
  wire  _T_91351; // @[OneHot.scala 66:30:@37128.4]
  wire  _T_91352; // @[OneHot.scala 66:30:@37129.4]
  wire  _T_91353; // @[OneHot.scala 66:30:@37130.4]
  wire  _T_91354; // @[OneHot.scala 66:30:@37131.4]
  wire  _T_91355; // @[OneHot.scala 66:30:@37132.4]
  wire  _T_91356; // @[OneHot.scala 66:30:@37133.4]
  wire  _T_91357; // @[OneHot.scala 66:30:@37134.4]
  wire [15:0] _T_91398; // @[Mux.scala 31:69:@37152.4]
  wire [15:0] _T_91399; // @[Mux.scala 31:69:@37153.4]
  wire [15:0] _T_91400; // @[Mux.scala 31:69:@37154.4]
  wire [15:0] _T_91401; // @[Mux.scala 31:69:@37155.4]
  wire [15:0] _T_91402; // @[Mux.scala 31:69:@37156.4]
  wire [15:0] _T_91403; // @[Mux.scala 31:69:@37157.4]
  wire [15:0] _T_91404; // @[Mux.scala 31:69:@37158.4]
  wire [15:0] _T_91405; // @[Mux.scala 31:69:@37159.4]
  wire [15:0] _T_91406; // @[Mux.scala 31:69:@37160.4]
  wire [15:0] _T_91407; // @[Mux.scala 31:69:@37161.4]
  wire [15:0] _T_91408; // @[Mux.scala 31:69:@37162.4]
  wire [15:0] _T_91409; // @[Mux.scala 31:69:@37163.4]
  wire [15:0] _T_91410; // @[Mux.scala 31:69:@37164.4]
  wire [15:0] _T_91411; // @[Mux.scala 31:69:@37165.4]
  wire [15:0] _T_91412; // @[Mux.scala 31:69:@37166.4]
  wire [15:0] _T_91413; // @[Mux.scala 31:69:@37167.4]
  wire  _T_91414; // @[OneHot.scala 66:30:@37168.4]
  wire  _T_91415; // @[OneHot.scala 66:30:@37169.4]
  wire  _T_91416; // @[OneHot.scala 66:30:@37170.4]
  wire  _T_91417; // @[OneHot.scala 66:30:@37171.4]
  wire  _T_91418; // @[OneHot.scala 66:30:@37172.4]
  wire  _T_91419; // @[OneHot.scala 66:30:@37173.4]
  wire  _T_91420; // @[OneHot.scala 66:30:@37174.4]
  wire  _T_91421; // @[OneHot.scala 66:30:@37175.4]
  wire  _T_91422; // @[OneHot.scala 66:30:@37176.4]
  wire  _T_91423; // @[OneHot.scala 66:30:@37177.4]
  wire  _T_91424; // @[OneHot.scala 66:30:@37178.4]
  wire  _T_91425; // @[OneHot.scala 66:30:@37179.4]
  wire  _T_91426; // @[OneHot.scala 66:30:@37180.4]
  wire  _T_91427; // @[OneHot.scala 66:30:@37181.4]
  wire  _T_91428; // @[OneHot.scala 66:30:@37182.4]
  wire  _T_91429; // @[OneHot.scala 66:30:@37183.4]
  wire [15:0] _T_91470; // @[Mux.scala 31:69:@37201.4]
  wire [15:0] _T_91471; // @[Mux.scala 31:69:@37202.4]
  wire [15:0] _T_91472; // @[Mux.scala 31:69:@37203.4]
  wire [15:0] _T_91473; // @[Mux.scala 31:69:@37204.4]
  wire [15:0] _T_91474; // @[Mux.scala 31:69:@37205.4]
  wire [15:0] _T_91475; // @[Mux.scala 31:69:@37206.4]
  wire [15:0] _T_91476; // @[Mux.scala 31:69:@37207.4]
  wire [15:0] _T_91477; // @[Mux.scala 31:69:@37208.4]
  wire [15:0] _T_91478; // @[Mux.scala 31:69:@37209.4]
  wire [15:0] _T_91479; // @[Mux.scala 31:69:@37210.4]
  wire [15:0] _T_91480; // @[Mux.scala 31:69:@37211.4]
  wire [15:0] _T_91481; // @[Mux.scala 31:69:@37212.4]
  wire [15:0] _T_91482; // @[Mux.scala 31:69:@37213.4]
  wire [15:0] _T_91483; // @[Mux.scala 31:69:@37214.4]
  wire [15:0] _T_91484; // @[Mux.scala 31:69:@37215.4]
  wire [15:0] _T_91485; // @[Mux.scala 31:69:@37216.4]
  wire  _T_91486; // @[OneHot.scala 66:30:@37217.4]
  wire  _T_91487; // @[OneHot.scala 66:30:@37218.4]
  wire  _T_91488; // @[OneHot.scala 66:30:@37219.4]
  wire  _T_91489; // @[OneHot.scala 66:30:@37220.4]
  wire  _T_91490; // @[OneHot.scala 66:30:@37221.4]
  wire  _T_91491; // @[OneHot.scala 66:30:@37222.4]
  wire  _T_91492; // @[OneHot.scala 66:30:@37223.4]
  wire  _T_91493; // @[OneHot.scala 66:30:@37224.4]
  wire  _T_91494; // @[OneHot.scala 66:30:@37225.4]
  wire  _T_91495; // @[OneHot.scala 66:30:@37226.4]
  wire  _T_91496; // @[OneHot.scala 66:30:@37227.4]
  wire  _T_91497; // @[OneHot.scala 66:30:@37228.4]
  wire  _T_91498; // @[OneHot.scala 66:30:@37229.4]
  wire  _T_91499; // @[OneHot.scala 66:30:@37230.4]
  wire  _T_91500; // @[OneHot.scala 66:30:@37231.4]
  wire  _T_91501; // @[OneHot.scala 66:30:@37232.4]
  wire [15:0] _T_91542; // @[Mux.scala 31:69:@37250.4]
  wire [15:0] _T_91543; // @[Mux.scala 31:69:@37251.4]
  wire [15:0] _T_91544; // @[Mux.scala 31:69:@37252.4]
  wire [15:0] _T_91545; // @[Mux.scala 31:69:@37253.4]
  wire [15:0] _T_91546; // @[Mux.scala 31:69:@37254.4]
  wire [15:0] _T_91547; // @[Mux.scala 31:69:@37255.4]
  wire [15:0] _T_91548; // @[Mux.scala 31:69:@37256.4]
  wire [15:0] _T_91549; // @[Mux.scala 31:69:@37257.4]
  wire [15:0] _T_91550; // @[Mux.scala 31:69:@37258.4]
  wire [15:0] _T_91551; // @[Mux.scala 31:69:@37259.4]
  wire [15:0] _T_91552; // @[Mux.scala 31:69:@37260.4]
  wire [15:0] _T_91553; // @[Mux.scala 31:69:@37261.4]
  wire [15:0] _T_91554; // @[Mux.scala 31:69:@37262.4]
  wire [15:0] _T_91555; // @[Mux.scala 31:69:@37263.4]
  wire [15:0] _T_91556; // @[Mux.scala 31:69:@37264.4]
  wire [15:0] _T_91557; // @[Mux.scala 31:69:@37265.4]
  wire  _T_91558; // @[OneHot.scala 66:30:@37266.4]
  wire  _T_91559; // @[OneHot.scala 66:30:@37267.4]
  wire  _T_91560; // @[OneHot.scala 66:30:@37268.4]
  wire  _T_91561; // @[OneHot.scala 66:30:@37269.4]
  wire  _T_91562; // @[OneHot.scala 66:30:@37270.4]
  wire  _T_91563; // @[OneHot.scala 66:30:@37271.4]
  wire  _T_91564; // @[OneHot.scala 66:30:@37272.4]
  wire  _T_91565; // @[OneHot.scala 66:30:@37273.4]
  wire  _T_91566; // @[OneHot.scala 66:30:@37274.4]
  wire  _T_91567; // @[OneHot.scala 66:30:@37275.4]
  wire  _T_91568; // @[OneHot.scala 66:30:@37276.4]
  wire  _T_91569; // @[OneHot.scala 66:30:@37277.4]
  wire  _T_91570; // @[OneHot.scala 66:30:@37278.4]
  wire  _T_91571; // @[OneHot.scala 66:30:@37279.4]
  wire  _T_91572; // @[OneHot.scala 66:30:@37280.4]
  wire  _T_91573; // @[OneHot.scala 66:30:@37281.4]
  wire [7:0] _T_91638; // @[Mux.scala 19:72:@37305.4]
  wire [15:0] _T_91646; // @[Mux.scala 19:72:@37313.4]
  wire [15:0] _T_91648; // @[Mux.scala 19:72:@37314.4]
  wire [7:0] _T_91655; // @[Mux.scala 19:72:@37321.4]
  wire [15:0] _T_91663; // @[Mux.scala 19:72:@37329.4]
  wire [15:0] _T_91665; // @[Mux.scala 19:72:@37330.4]
  wire [7:0] _T_91672; // @[Mux.scala 19:72:@37337.4]
  wire [15:0] _T_91680; // @[Mux.scala 19:72:@37345.4]
  wire [15:0] _T_91682; // @[Mux.scala 19:72:@37346.4]
  wire [7:0] _T_91689; // @[Mux.scala 19:72:@37353.4]
  wire [15:0] _T_91697; // @[Mux.scala 19:72:@37361.4]
  wire [15:0] _T_91699; // @[Mux.scala 19:72:@37362.4]
  wire [7:0] _T_91706; // @[Mux.scala 19:72:@37369.4]
  wire [15:0] _T_91714; // @[Mux.scala 19:72:@37377.4]
  wire [15:0] _T_91716; // @[Mux.scala 19:72:@37378.4]
  wire [7:0] _T_91723; // @[Mux.scala 19:72:@37385.4]
  wire [15:0] _T_91731; // @[Mux.scala 19:72:@37393.4]
  wire [15:0] _T_91733; // @[Mux.scala 19:72:@37394.4]
  wire [7:0] _T_91740; // @[Mux.scala 19:72:@37401.4]
  wire [15:0] _T_91748; // @[Mux.scala 19:72:@37409.4]
  wire [15:0] _T_91750; // @[Mux.scala 19:72:@37410.4]
  wire [7:0] _T_91757; // @[Mux.scala 19:72:@37417.4]
  wire [15:0] _T_91765; // @[Mux.scala 19:72:@37425.4]
  wire [15:0] _T_91767; // @[Mux.scala 19:72:@37426.4]
  wire [7:0] _T_91774; // @[Mux.scala 19:72:@37433.4]
  wire [15:0] _T_91782; // @[Mux.scala 19:72:@37441.4]
  wire [15:0] _T_91784; // @[Mux.scala 19:72:@37442.4]
  wire [7:0] _T_91791; // @[Mux.scala 19:72:@37449.4]
  wire [15:0] _T_91799; // @[Mux.scala 19:72:@37457.4]
  wire [15:0] _T_91801; // @[Mux.scala 19:72:@37458.4]
  wire [7:0] _T_91808; // @[Mux.scala 19:72:@37465.4]
  wire [15:0] _T_91816; // @[Mux.scala 19:72:@37473.4]
  wire [15:0] _T_91818; // @[Mux.scala 19:72:@37474.4]
  wire [7:0] _T_91825; // @[Mux.scala 19:72:@37481.4]
  wire [15:0] _T_91833; // @[Mux.scala 19:72:@37489.4]
  wire [15:0] _T_91835; // @[Mux.scala 19:72:@37490.4]
  wire [7:0] _T_91842; // @[Mux.scala 19:72:@37497.4]
  wire [15:0] _T_91850; // @[Mux.scala 19:72:@37505.4]
  wire [15:0] _T_91852; // @[Mux.scala 19:72:@37506.4]
  wire [7:0] _T_91859; // @[Mux.scala 19:72:@37513.4]
  wire [15:0] _T_91867; // @[Mux.scala 19:72:@37521.4]
  wire [15:0] _T_91869; // @[Mux.scala 19:72:@37522.4]
  wire [7:0] _T_91876; // @[Mux.scala 19:72:@37529.4]
  wire [15:0] _T_91884; // @[Mux.scala 19:72:@37537.4]
  wire [15:0] _T_91886; // @[Mux.scala 19:72:@37538.4]
  wire [7:0] _T_91893; // @[Mux.scala 19:72:@37545.4]
  wire [15:0] _T_91901; // @[Mux.scala 19:72:@37553.4]
  wire [15:0] _T_91903; // @[Mux.scala 19:72:@37554.4]
  wire [15:0] _T_91904; // @[Mux.scala 19:72:@37555.4]
  wire [15:0] _T_91905; // @[Mux.scala 19:72:@37556.4]
  wire [15:0] _T_91906; // @[Mux.scala 19:72:@37557.4]
  wire [15:0] _T_91907; // @[Mux.scala 19:72:@37558.4]
  wire [15:0] _T_91908; // @[Mux.scala 19:72:@37559.4]
  wire [15:0] _T_91909; // @[Mux.scala 19:72:@37560.4]
  wire [15:0] _T_91910; // @[Mux.scala 19:72:@37561.4]
  wire [15:0] _T_91911; // @[Mux.scala 19:72:@37562.4]
  wire [15:0] _T_91912; // @[Mux.scala 19:72:@37563.4]
  wire [15:0] _T_91913; // @[Mux.scala 19:72:@37564.4]
  wire [15:0] _T_91914; // @[Mux.scala 19:72:@37565.4]
  wire [15:0] _T_91915; // @[Mux.scala 19:72:@37566.4]
  wire [15:0] _T_91916; // @[Mux.scala 19:72:@37567.4]
  wire [15:0] _T_91917; // @[Mux.scala 19:72:@37568.4]
  wire [15:0] _T_91918; // @[Mux.scala 19:72:@37569.4]
  wire  priorityLoadRequest_0; // @[Mux.scala 19:72:@37573.4]
  wire  priorityLoadRequest_1; // @[Mux.scala 19:72:@37575.4]
  wire  priorityLoadRequest_2; // @[Mux.scala 19:72:@37577.4]
  wire  priorityLoadRequest_3; // @[Mux.scala 19:72:@37579.4]
  wire  priorityLoadRequest_4; // @[Mux.scala 19:72:@37581.4]
  wire  priorityLoadRequest_5; // @[Mux.scala 19:72:@37583.4]
  wire  priorityLoadRequest_6; // @[Mux.scala 19:72:@37585.4]
  wire  priorityLoadRequest_7; // @[Mux.scala 19:72:@37587.4]
  wire  priorityLoadRequest_8; // @[Mux.scala 19:72:@37589.4]
  wire  priorityLoadRequest_9; // @[Mux.scala 19:72:@37591.4]
  wire  priorityLoadRequest_10; // @[Mux.scala 19:72:@37593.4]
  wire  priorityLoadRequest_11; // @[Mux.scala 19:72:@37595.4]
  wire  priorityLoadRequest_12; // @[Mux.scala 19:72:@37597.4]
  wire  priorityLoadRequest_13; // @[Mux.scala 19:72:@37599.4]
  wire  priorityLoadRequest_14; // @[Mux.scala 19:72:@37601.4]
  wire  priorityLoadRequest_15; // @[Mux.scala 19:72:@37603.4]
  wire  _T_92186; // @[AxiLoadQueue.scala 212:39:@37627.6]
  wire  _GEN_1920; // @[AxiLoadQueue.scala 212:70:@37628.6]
  wire  _GEN_1921; // @[AxiLoadQueue.scala 210:22:@37623.4]
  wire  _T_92189; // @[AxiLoadQueue.scala 212:39:@37635.6]
  wire  _GEN_1922; // @[AxiLoadQueue.scala 212:70:@37636.6]
  wire  _GEN_1923; // @[AxiLoadQueue.scala 210:22:@37631.4]
  wire  _T_92192; // @[AxiLoadQueue.scala 212:39:@37643.6]
  wire  _GEN_1924; // @[AxiLoadQueue.scala 212:70:@37644.6]
  wire  _GEN_1925; // @[AxiLoadQueue.scala 210:22:@37639.4]
  wire  _T_92195; // @[AxiLoadQueue.scala 212:39:@37651.6]
  wire  _GEN_1926; // @[AxiLoadQueue.scala 212:70:@37652.6]
  wire  _GEN_1927; // @[AxiLoadQueue.scala 210:22:@37647.4]
  wire  _T_92198; // @[AxiLoadQueue.scala 212:39:@37659.6]
  wire  _GEN_1928; // @[AxiLoadQueue.scala 212:70:@37660.6]
  wire  _GEN_1929; // @[AxiLoadQueue.scala 210:22:@37655.4]
  wire  _T_92201; // @[AxiLoadQueue.scala 212:39:@37667.6]
  wire  _GEN_1930; // @[AxiLoadQueue.scala 212:70:@37668.6]
  wire  _GEN_1931; // @[AxiLoadQueue.scala 210:22:@37663.4]
  wire  _T_92204; // @[AxiLoadQueue.scala 212:39:@37675.6]
  wire  _GEN_1932; // @[AxiLoadQueue.scala 212:70:@37676.6]
  wire  _GEN_1933; // @[AxiLoadQueue.scala 210:22:@37671.4]
  wire  _T_92207; // @[AxiLoadQueue.scala 212:39:@37683.6]
  wire  _GEN_1934; // @[AxiLoadQueue.scala 212:70:@37684.6]
  wire  _GEN_1935; // @[AxiLoadQueue.scala 210:22:@37679.4]
  wire  _T_92210; // @[AxiLoadQueue.scala 212:39:@37691.6]
  wire  _GEN_1936; // @[AxiLoadQueue.scala 212:70:@37692.6]
  wire  _GEN_1937; // @[AxiLoadQueue.scala 210:22:@37687.4]
  wire  _T_92213; // @[AxiLoadQueue.scala 212:39:@37699.6]
  wire  _GEN_1938; // @[AxiLoadQueue.scala 212:70:@37700.6]
  wire  _GEN_1939; // @[AxiLoadQueue.scala 210:22:@37695.4]
  wire  _T_92216; // @[AxiLoadQueue.scala 212:39:@37707.6]
  wire  _GEN_1940; // @[AxiLoadQueue.scala 212:70:@37708.6]
  wire  _GEN_1941; // @[AxiLoadQueue.scala 210:22:@37703.4]
  wire  _T_92219; // @[AxiLoadQueue.scala 212:39:@37715.6]
  wire  _GEN_1942; // @[AxiLoadQueue.scala 212:70:@37716.6]
  wire  _GEN_1943; // @[AxiLoadQueue.scala 210:22:@37711.4]
  wire  _T_92222; // @[AxiLoadQueue.scala 212:39:@37723.6]
  wire  _GEN_1944; // @[AxiLoadQueue.scala 212:70:@37724.6]
  wire  _GEN_1945; // @[AxiLoadQueue.scala 210:22:@37719.4]
  wire  _T_92225; // @[AxiLoadQueue.scala 212:39:@37731.6]
  wire  _GEN_1946; // @[AxiLoadQueue.scala 212:70:@37732.6]
  wire  _GEN_1947; // @[AxiLoadQueue.scala 210:22:@37727.4]
  wire  _T_92228; // @[AxiLoadQueue.scala 212:39:@37739.6]
  wire  _GEN_1948; // @[AxiLoadQueue.scala 212:70:@37740.6]
  wire  _GEN_1949; // @[AxiLoadQueue.scala 210:22:@37735.4]
  wire  _T_92231; // @[AxiLoadQueue.scala 212:39:@37747.6]
  wire  _GEN_1950; // @[AxiLoadQueue.scala 212:70:@37748.6]
  wire  _GEN_1951; // @[AxiLoadQueue.scala 210:22:@37743.4]
  wire [3:0] _T_92249; // @[Mux.scala 31:69:@37751.4]
  wire [3:0] _T_92250; // @[Mux.scala 31:69:@37752.4]
  wire [3:0] _T_92251; // @[Mux.scala 31:69:@37753.4]
  wire [3:0] _T_92252; // @[Mux.scala 31:69:@37754.4]
  wire [3:0] _T_92253; // @[Mux.scala 31:69:@37755.4]
  wire [3:0] _T_92254; // @[Mux.scala 31:69:@37756.4]
  wire [3:0] _T_92255; // @[Mux.scala 31:69:@37757.4]
  wire [3:0] _T_92256; // @[Mux.scala 31:69:@37758.4]
  wire [3:0] _T_92257; // @[Mux.scala 31:69:@37759.4]
  wire [3:0] _T_92258; // @[Mux.scala 31:69:@37760.4]
  wire [3:0] _T_92259; // @[Mux.scala 31:69:@37761.4]
  wire [3:0] _T_92260; // @[Mux.scala 31:69:@37762.4]
  wire [3:0] _T_92261; // @[Mux.scala 31:69:@37763.4]
  wire [3:0] _T_92262; // @[Mux.scala 31:69:@37764.4]
  wire [3:0] _T_92263; // @[Mux.scala 31:69:@37765.4]
  wire  _T_92266; // @[AxiLoadQueue.scala 222:60:@37768.4]
  wire  _T_92267; // @[AxiLoadQueue.scala 222:60:@37769.4]
  wire  _T_92268; // @[AxiLoadQueue.scala 222:60:@37770.4]
  wire  _T_92269; // @[AxiLoadQueue.scala 222:60:@37771.4]
  wire  _T_92270; // @[AxiLoadQueue.scala 222:60:@37772.4]
  wire  _T_92271; // @[AxiLoadQueue.scala 222:60:@37773.4]
  wire  _T_92272; // @[AxiLoadQueue.scala 222:60:@37774.4]
  wire  _T_92273; // @[AxiLoadQueue.scala 222:60:@37775.4]
  wire  _T_92274; // @[AxiLoadQueue.scala 222:60:@37776.4]
  wire  _T_92275; // @[AxiLoadQueue.scala 222:60:@37777.4]
  wire  _T_92276; // @[AxiLoadQueue.scala 222:60:@37778.4]
  wire  _T_92277; // @[AxiLoadQueue.scala 222:60:@37779.4]
  wire  _T_92278; // @[AxiLoadQueue.scala 222:60:@37780.4]
  wire  _T_92279; // @[AxiLoadQueue.scala 222:60:@37781.4]
  wire [30:0] _GEN_1953; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1954; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1955; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1956; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1957; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1958; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1959; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1960; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1961; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1962; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1963; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1964; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1965; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [30:0] _GEN_1966; // @[AxiLoadQueue.scala 223:20:@37799.4]
  wire [7:0] _T_92405; // @[AxiLoadQueue.scala 251:58:@37965.8]
  wire [15:0] _T_92413; // @[AxiLoadQueue.scala 251:58:@37973.8]
  wire [7:0] _T_92420; // @[AxiLoadQueue.scala 251:96:@37980.8]
  wire [15:0] _T_92428; // @[AxiLoadQueue.scala 251:96:@37988.8]
  wire  _T_92429; // @[AxiLoadQueue.scala 251:61:@37989.8]
  wire  _T_92430; // @[AxiLoadQueue.scala 250:64:@37990.8]
  wire  _GEN_2001; // @[AxiLoadQueue.scala 243:104:@37922.6]
  wire  bypassRequest_0; // @[AxiLoadQueue.scala 242:71:@37916.4]
  wire  _GEN_1968; // @[AxiLoadQueue.scala 230:34:@37804.6]
  wire  _GEN_1969; // @[AxiLoadQueue.scala 228:23:@37800.4]
  wire [7:0] _T_92489; // @[AxiLoadQueue.scala 251:58:@38047.8]
  wire [15:0] _T_92497; // @[AxiLoadQueue.scala 251:58:@38055.8]
  wire [7:0] _T_92504; // @[AxiLoadQueue.scala 251:96:@38062.8]
  wire [15:0] _T_92512; // @[AxiLoadQueue.scala 251:96:@38070.8]
  wire  _T_92513; // @[AxiLoadQueue.scala 251:61:@38071.8]
  wire  _T_92514; // @[AxiLoadQueue.scala 250:64:@38072.8]
  wire  _GEN_2005; // @[AxiLoadQueue.scala 243:104:@38004.6]
  wire  bypassRequest_1; // @[AxiLoadQueue.scala 242:71:@37998.4]
  wire  _GEN_1970; // @[AxiLoadQueue.scala 230:34:@37811.6]
  wire  _GEN_1971; // @[AxiLoadQueue.scala 228:23:@37807.4]
  wire [7:0] _T_92573; // @[AxiLoadQueue.scala 251:58:@38129.8]
  wire [15:0] _T_92581; // @[AxiLoadQueue.scala 251:58:@38137.8]
  wire [7:0] _T_92588; // @[AxiLoadQueue.scala 251:96:@38144.8]
  wire [15:0] _T_92596; // @[AxiLoadQueue.scala 251:96:@38152.8]
  wire  _T_92597; // @[AxiLoadQueue.scala 251:61:@38153.8]
  wire  _T_92598; // @[AxiLoadQueue.scala 250:64:@38154.8]
  wire  _GEN_2009; // @[AxiLoadQueue.scala 243:104:@38086.6]
  wire  bypassRequest_2; // @[AxiLoadQueue.scala 242:71:@38080.4]
  wire  _GEN_1972; // @[AxiLoadQueue.scala 230:34:@37818.6]
  wire  _GEN_1973; // @[AxiLoadQueue.scala 228:23:@37814.4]
  wire [7:0] _T_92657; // @[AxiLoadQueue.scala 251:58:@38211.8]
  wire [15:0] _T_92665; // @[AxiLoadQueue.scala 251:58:@38219.8]
  wire [7:0] _T_92672; // @[AxiLoadQueue.scala 251:96:@38226.8]
  wire [15:0] _T_92680; // @[AxiLoadQueue.scala 251:96:@38234.8]
  wire  _T_92681; // @[AxiLoadQueue.scala 251:61:@38235.8]
  wire  _T_92682; // @[AxiLoadQueue.scala 250:64:@38236.8]
  wire  _GEN_2013; // @[AxiLoadQueue.scala 243:104:@38168.6]
  wire  bypassRequest_3; // @[AxiLoadQueue.scala 242:71:@38162.4]
  wire  _GEN_1974; // @[AxiLoadQueue.scala 230:34:@37825.6]
  wire  _GEN_1975; // @[AxiLoadQueue.scala 228:23:@37821.4]
  wire [7:0] _T_92741; // @[AxiLoadQueue.scala 251:58:@38293.8]
  wire [15:0] _T_92749; // @[AxiLoadQueue.scala 251:58:@38301.8]
  wire [7:0] _T_92756; // @[AxiLoadQueue.scala 251:96:@38308.8]
  wire [15:0] _T_92764; // @[AxiLoadQueue.scala 251:96:@38316.8]
  wire  _T_92765; // @[AxiLoadQueue.scala 251:61:@38317.8]
  wire  _T_92766; // @[AxiLoadQueue.scala 250:64:@38318.8]
  wire  _GEN_2017; // @[AxiLoadQueue.scala 243:104:@38250.6]
  wire  bypassRequest_4; // @[AxiLoadQueue.scala 242:71:@38244.4]
  wire  _GEN_1976; // @[AxiLoadQueue.scala 230:34:@37832.6]
  wire  _GEN_1977; // @[AxiLoadQueue.scala 228:23:@37828.4]
  wire [7:0] _T_92825; // @[AxiLoadQueue.scala 251:58:@38375.8]
  wire [15:0] _T_92833; // @[AxiLoadQueue.scala 251:58:@38383.8]
  wire [7:0] _T_92840; // @[AxiLoadQueue.scala 251:96:@38390.8]
  wire [15:0] _T_92848; // @[AxiLoadQueue.scala 251:96:@38398.8]
  wire  _T_92849; // @[AxiLoadQueue.scala 251:61:@38399.8]
  wire  _T_92850; // @[AxiLoadQueue.scala 250:64:@38400.8]
  wire  _GEN_2021; // @[AxiLoadQueue.scala 243:104:@38332.6]
  wire  bypassRequest_5; // @[AxiLoadQueue.scala 242:71:@38326.4]
  wire  _GEN_1978; // @[AxiLoadQueue.scala 230:34:@37839.6]
  wire  _GEN_1979; // @[AxiLoadQueue.scala 228:23:@37835.4]
  wire [7:0] _T_92909; // @[AxiLoadQueue.scala 251:58:@38457.8]
  wire [15:0] _T_92917; // @[AxiLoadQueue.scala 251:58:@38465.8]
  wire [7:0] _T_92924; // @[AxiLoadQueue.scala 251:96:@38472.8]
  wire [15:0] _T_92932; // @[AxiLoadQueue.scala 251:96:@38480.8]
  wire  _T_92933; // @[AxiLoadQueue.scala 251:61:@38481.8]
  wire  _T_92934; // @[AxiLoadQueue.scala 250:64:@38482.8]
  wire  _GEN_2025; // @[AxiLoadQueue.scala 243:104:@38414.6]
  wire  bypassRequest_6; // @[AxiLoadQueue.scala 242:71:@38408.4]
  wire  _GEN_1980; // @[AxiLoadQueue.scala 230:34:@37846.6]
  wire  _GEN_1981; // @[AxiLoadQueue.scala 228:23:@37842.4]
  wire [7:0] _T_92993; // @[AxiLoadQueue.scala 251:58:@38539.8]
  wire [15:0] _T_93001; // @[AxiLoadQueue.scala 251:58:@38547.8]
  wire [7:0] _T_93008; // @[AxiLoadQueue.scala 251:96:@38554.8]
  wire [15:0] _T_93016; // @[AxiLoadQueue.scala 251:96:@38562.8]
  wire  _T_93017; // @[AxiLoadQueue.scala 251:61:@38563.8]
  wire  _T_93018; // @[AxiLoadQueue.scala 250:64:@38564.8]
  wire  _GEN_2029; // @[AxiLoadQueue.scala 243:104:@38496.6]
  wire  bypassRequest_7; // @[AxiLoadQueue.scala 242:71:@38490.4]
  wire  _GEN_1982; // @[AxiLoadQueue.scala 230:34:@37853.6]
  wire  _GEN_1983; // @[AxiLoadQueue.scala 228:23:@37849.4]
  wire [7:0] _T_93077; // @[AxiLoadQueue.scala 251:58:@38621.8]
  wire [15:0] _T_93085; // @[AxiLoadQueue.scala 251:58:@38629.8]
  wire [7:0] _T_93092; // @[AxiLoadQueue.scala 251:96:@38636.8]
  wire [15:0] _T_93100; // @[AxiLoadQueue.scala 251:96:@38644.8]
  wire  _T_93101; // @[AxiLoadQueue.scala 251:61:@38645.8]
  wire  _T_93102; // @[AxiLoadQueue.scala 250:64:@38646.8]
  wire  _GEN_2033; // @[AxiLoadQueue.scala 243:104:@38578.6]
  wire  bypassRequest_8; // @[AxiLoadQueue.scala 242:71:@38572.4]
  wire  _GEN_1984; // @[AxiLoadQueue.scala 230:34:@37860.6]
  wire  _GEN_1985; // @[AxiLoadQueue.scala 228:23:@37856.4]
  wire [7:0] _T_93161; // @[AxiLoadQueue.scala 251:58:@38703.8]
  wire [15:0] _T_93169; // @[AxiLoadQueue.scala 251:58:@38711.8]
  wire [7:0] _T_93176; // @[AxiLoadQueue.scala 251:96:@38718.8]
  wire [15:0] _T_93184; // @[AxiLoadQueue.scala 251:96:@38726.8]
  wire  _T_93185; // @[AxiLoadQueue.scala 251:61:@38727.8]
  wire  _T_93186; // @[AxiLoadQueue.scala 250:64:@38728.8]
  wire  _GEN_2037; // @[AxiLoadQueue.scala 243:104:@38660.6]
  wire  bypassRequest_9; // @[AxiLoadQueue.scala 242:71:@38654.4]
  wire  _GEN_1986; // @[AxiLoadQueue.scala 230:34:@37867.6]
  wire  _GEN_1987; // @[AxiLoadQueue.scala 228:23:@37863.4]
  wire [7:0] _T_93245; // @[AxiLoadQueue.scala 251:58:@38785.8]
  wire [15:0] _T_93253; // @[AxiLoadQueue.scala 251:58:@38793.8]
  wire [7:0] _T_93260; // @[AxiLoadQueue.scala 251:96:@38800.8]
  wire [15:0] _T_93268; // @[AxiLoadQueue.scala 251:96:@38808.8]
  wire  _T_93269; // @[AxiLoadQueue.scala 251:61:@38809.8]
  wire  _T_93270; // @[AxiLoadQueue.scala 250:64:@38810.8]
  wire  _GEN_2041; // @[AxiLoadQueue.scala 243:104:@38742.6]
  wire  bypassRequest_10; // @[AxiLoadQueue.scala 242:71:@38736.4]
  wire  _GEN_1988; // @[AxiLoadQueue.scala 230:34:@37874.6]
  wire  _GEN_1989; // @[AxiLoadQueue.scala 228:23:@37870.4]
  wire [7:0] _T_93329; // @[AxiLoadQueue.scala 251:58:@38867.8]
  wire [15:0] _T_93337; // @[AxiLoadQueue.scala 251:58:@38875.8]
  wire [7:0] _T_93344; // @[AxiLoadQueue.scala 251:96:@38882.8]
  wire [15:0] _T_93352; // @[AxiLoadQueue.scala 251:96:@38890.8]
  wire  _T_93353; // @[AxiLoadQueue.scala 251:61:@38891.8]
  wire  _T_93354; // @[AxiLoadQueue.scala 250:64:@38892.8]
  wire  _GEN_2045; // @[AxiLoadQueue.scala 243:104:@38824.6]
  wire  bypassRequest_11; // @[AxiLoadQueue.scala 242:71:@38818.4]
  wire  _GEN_1990; // @[AxiLoadQueue.scala 230:34:@37881.6]
  wire  _GEN_1991; // @[AxiLoadQueue.scala 228:23:@37877.4]
  wire [7:0] _T_93413; // @[AxiLoadQueue.scala 251:58:@38949.8]
  wire [15:0] _T_93421; // @[AxiLoadQueue.scala 251:58:@38957.8]
  wire [7:0] _T_93428; // @[AxiLoadQueue.scala 251:96:@38964.8]
  wire [15:0] _T_93436; // @[AxiLoadQueue.scala 251:96:@38972.8]
  wire  _T_93437; // @[AxiLoadQueue.scala 251:61:@38973.8]
  wire  _T_93438; // @[AxiLoadQueue.scala 250:64:@38974.8]
  wire  _GEN_2049; // @[AxiLoadQueue.scala 243:104:@38906.6]
  wire  bypassRequest_12; // @[AxiLoadQueue.scala 242:71:@38900.4]
  wire  _GEN_1992; // @[AxiLoadQueue.scala 230:34:@37888.6]
  wire  _GEN_1993; // @[AxiLoadQueue.scala 228:23:@37884.4]
  wire [7:0] _T_93497; // @[AxiLoadQueue.scala 251:58:@39031.8]
  wire [15:0] _T_93505; // @[AxiLoadQueue.scala 251:58:@39039.8]
  wire [7:0] _T_93512; // @[AxiLoadQueue.scala 251:96:@39046.8]
  wire [15:0] _T_93520; // @[AxiLoadQueue.scala 251:96:@39054.8]
  wire  _T_93521; // @[AxiLoadQueue.scala 251:61:@39055.8]
  wire  _T_93522; // @[AxiLoadQueue.scala 250:64:@39056.8]
  wire  _GEN_2053; // @[AxiLoadQueue.scala 243:104:@38988.6]
  wire  bypassRequest_13; // @[AxiLoadQueue.scala 242:71:@38982.4]
  wire  _GEN_1994; // @[AxiLoadQueue.scala 230:34:@37895.6]
  wire  _GEN_1995; // @[AxiLoadQueue.scala 228:23:@37891.4]
  wire [7:0] _T_93581; // @[AxiLoadQueue.scala 251:58:@39113.8]
  wire [15:0] _T_93589; // @[AxiLoadQueue.scala 251:58:@39121.8]
  wire [7:0] _T_93596; // @[AxiLoadQueue.scala 251:96:@39128.8]
  wire [15:0] _T_93604; // @[AxiLoadQueue.scala 251:96:@39136.8]
  wire  _T_93605; // @[AxiLoadQueue.scala 251:61:@39137.8]
  wire  _T_93606; // @[AxiLoadQueue.scala 250:64:@39138.8]
  wire  _GEN_2057; // @[AxiLoadQueue.scala 243:104:@39070.6]
  wire  bypassRequest_14; // @[AxiLoadQueue.scala 242:71:@39064.4]
  wire  _GEN_1996; // @[AxiLoadQueue.scala 230:34:@37902.6]
  wire  _GEN_1997; // @[AxiLoadQueue.scala 228:23:@37898.4]
  wire [7:0] _T_93665; // @[AxiLoadQueue.scala 251:58:@39195.8]
  wire [15:0] _T_93673; // @[AxiLoadQueue.scala 251:58:@39203.8]
  wire [7:0] _T_93680; // @[AxiLoadQueue.scala 251:96:@39210.8]
  wire [15:0] _T_93688; // @[AxiLoadQueue.scala 251:96:@39218.8]
  wire  _T_93689; // @[AxiLoadQueue.scala 251:61:@39219.8]
  wire  _T_93690; // @[AxiLoadQueue.scala 250:64:@39220.8]
  wire  _GEN_2061; // @[AxiLoadQueue.scala 243:104:@39152.6]
  wire  bypassRequest_15; // @[AxiLoadQueue.scala 242:71:@39146.4]
  wire  _GEN_1998; // @[AxiLoadQueue.scala 230:34:@37909.6]
  wire  _GEN_1999; // @[AxiLoadQueue.scala 228:23:@37905.4]
  wire  _T_93693; // @[AxiLoadQueue.scala 262:69:@39228.6]
  wire  _T_93694; // @[AxiLoadQueue.scala 262:45:@39229.6]
  wire  _T_93695; // @[AxiLoadQueue.scala 262:78:@39230.6]
  wire  _GEN_2064; // @[AxiLoadQueue.scala 262:99:@39231.6]
  wire  _GEN_2065; // @[AxiLoadQueue.scala 260:25:@39224.4]
  wire  _T_93699; // @[AxiLoadQueue.scala 262:69:@39238.6]
  wire  _T_93700; // @[AxiLoadQueue.scala 262:45:@39239.6]
  wire  _T_93701; // @[AxiLoadQueue.scala 262:78:@39240.6]
  wire  _GEN_2066; // @[AxiLoadQueue.scala 262:99:@39241.6]
  wire  _GEN_2067; // @[AxiLoadQueue.scala 260:25:@39234.4]
  wire  _T_93705; // @[AxiLoadQueue.scala 262:69:@39248.6]
  wire  _T_93706; // @[AxiLoadQueue.scala 262:45:@39249.6]
  wire  _T_93707; // @[AxiLoadQueue.scala 262:78:@39250.6]
  wire  _GEN_2068; // @[AxiLoadQueue.scala 262:99:@39251.6]
  wire  _GEN_2069; // @[AxiLoadQueue.scala 260:25:@39244.4]
  wire  _T_93711; // @[AxiLoadQueue.scala 262:69:@39258.6]
  wire  _T_93712; // @[AxiLoadQueue.scala 262:45:@39259.6]
  wire  _T_93713; // @[AxiLoadQueue.scala 262:78:@39260.6]
  wire  _GEN_2070; // @[AxiLoadQueue.scala 262:99:@39261.6]
  wire  _GEN_2071; // @[AxiLoadQueue.scala 260:25:@39254.4]
  wire  _T_93717; // @[AxiLoadQueue.scala 262:69:@39268.6]
  wire  _T_93718; // @[AxiLoadQueue.scala 262:45:@39269.6]
  wire  _T_93719; // @[AxiLoadQueue.scala 262:78:@39270.6]
  wire  _GEN_2072; // @[AxiLoadQueue.scala 262:99:@39271.6]
  wire  _GEN_2073; // @[AxiLoadQueue.scala 260:25:@39264.4]
  wire  _T_93723; // @[AxiLoadQueue.scala 262:69:@39278.6]
  wire  _T_93724; // @[AxiLoadQueue.scala 262:45:@39279.6]
  wire  _T_93725; // @[AxiLoadQueue.scala 262:78:@39280.6]
  wire  _GEN_2074; // @[AxiLoadQueue.scala 262:99:@39281.6]
  wire  _GEN_2075; // @[AxiLoadQueue.scala 260:25:@39274.4]
  wire  _T_93729; // @[AxiLoadQueue.scala 262:69:@39288.6]
  wire  _T_93730; // @[AxiLoadQueue.scala 262:45:@39289.6]
  wire  _T_93731; // @[AxiLoadQueue.scala 262:78:@39290.6]
  wire  _GEN_2076; // @[AxiLoadQueue.scala 262:99:@39291.6]
  wire  _GEN_2077; // @[AxiLoadQueue.scala 260:25:@39284.4]
  wire  _T_93735; // @[AxiLoadQueue.scala 262:69:@39298.6]
  wire  _T_93736; // @[AxiLoadQueue.scala 262:45:@39299.6]
  wire  _T_93737; // @[AxiLoadQueue.scala 262:78:@39300.6]
  wire  _GEN_2078; // @[AxiLoadQueue.scala 262:99:@39301.6]
  wire  _GEN_2079; // @[AxiLoadQueue.scala 260:25:@39294.4]
  wire  _T_93741; // @[AxiLoadQueue.scala 262:69:@39308.6]
  wire  _T_93742; // @[AxiLoadQueue.scala 262:45:@39309.6]
  wire  _T_93743; // @[AxiLoadQueue.scala 262:78:@39310.6]
  wire  _GEN_2080; // @[AxiLoadQueue.scala 262:99:@39311.6]
  wire  _GEN_2081; // @[AxiLoadQueue.scala 260:25:@39304.4]
  wire  _T_93747; // @[AxiLoadQueue.scala 262:69:@39318.6]
  wire  _T_93748; // @[AxiLoadQueue.scala 262:45:@39319.6]
  wire  _T_93749; // @[AxiLoadQueue.scala 262:78:@39320.6]
  wire  _GEN_2082; // @[AxiLoadQueue.scala 262:99:@39321.6]
  wire  _GEN_2083; // @[AxiLoadQueue.scala 260:25:@39314.4]
  wire  _T_93753; // @[AxiLoadQueue.scala 262:69:@39328.6]
  wire  _T_93754; // @[AxiLoadQueue.scala 262:45:@39329.6]
  wire  _T_93755; // @[AxiLoadQueue.scala 262:78:@39330.6]
  wire  _GEN_2084; // @[AxiLoadQueue.scala 262:99:@39331.6]
  wire  _GEN_2085; // @[AxiLoadQueue.scala 260:25:@39324.4]
  wire  _T_93759; // @[AxiLoadQueue.scala 262:69:@39338.6]
  wire  _T_93760; // @[AxiLoadQueue.scala 262:45:@39339.6]
  wire  _T_93761; // @[AxiLoadQueue.scala 262:78:@39340.6]
  wire  _GEN_2086; // @[AxiLoadQueue.scala 262:99:@39341.6]
  wire  _GEN_2087; // @[AxiLoadQueue.scala 260:25:@39334.4]
  wire  _T_93765; // @[AxiLoadQueue.scala 262:69:@39348.6]
  wire  _T_93766; // @[AxiLoadQueue.scala 262:45:@39349.6]
  wire  _T_93767; // @[AxiLoadQueue.scala 262:78:@39350.6]
  wire  _GEN_2088; // @[AxiLoadQueue.scala 262:99:@39351.6]
  wire  _GEN_2089; // @[AxiLoadQueue.scala 260:25:@39344.4]
  wire  _T_93771; // @[AxiLoadQueue.scala 262:69:@39358.6]
  wire  _T_93772; // @[AxiLoadQueue.scala 262:45:@39359.6]
  wire  _T_93773; // @[AxiLoadQueue.scala 262:78:@39360.6]
  wire  _GEN_2090; // @[AxiLoadQueue.scala 262:99:@39361.6]
  wire  _GEN_2091; // @[AxiLoadQueue.scala 260:25:@39354.4]
  wire  _T_93777; // @[AxiLoadQueue.scala 262:69:@39368.6]
  wire  _T_93778; // @[AxiLoadQueue.scala 262:45:@39369.6]
  wire  _T_93779; // @[AxiLoadQueue.scala 262:78:@39370.6]
  wire  _GEN_2092; // @[AxiLoadQueue.scala 262:99:@39371.6]
  wire  _GEN_2093; // @[AxiLoadQueue.scala 260:25:@39364.4]
  wire  _T_93783; // @[AxiLoadQueue.scala 262:69:@39378.6]
  wire  _T_93784; // @[AxiLoadQueue.scala 262:45:@39379.6]
  wire  _T_93785; // @[AxiLoadQueue.scala 262:78:@39380.6]
  wire  _GEN_2094; // @[AxiLoadQueue.scala 262:99:@39381.6]
  wire  _GEN_2095; // @[AxiLoadQueue.scala 260:25:@39374.4]
  wire [31:0] _GEN_2096; // @[AxiLoadQueue.scala 270:79:@39390.6]
  wire [31:0] _GEN_2097; // @[AxiLoadQueue.scala 268:32:@39384.4]
  wire [31:0] _GEN_2098; // @[AxiLoadQueue.scala 270:79:@39399.6]
  wire [31:0] _GEN_2099; // @[AxiLoadQueue.scala 268:32:@39393.4]
  wire [31:0] _GEN_2100; // @[AxiLoadQueue.scala 270:79:@39408.6]
  wire [31:0] _GEN_2101; // @[AxiLoadQueue.scala 268:32:@39402.4]
  wire [31:0] _GEN_2102; // @[AxiLoadQueue.scala 270:79:@39417.6]
  wire [31:0] _GEN_2103; // @[AxiLoadQueue.scala 268:32:@39411.4]
  wire [31:0] _GEN_2104; // @[AxiLoadQueue.scala 270:79:@39426.6]
  wire [31:0] _GEN_2105; // @[AxiLoadQueue.scala 268:32:@39420.4]
  wire [31:0] _GEN_2106; // @[AxiLoadQueue.scala 270:79:@39435.6]
  wire [31:0] _GEN_2107; // @[AxiLoadQueue.scala 268:32:@39429.4]
  wire [31:0] _GEN_2108; // @[AxiLoadQueue.scala 270:79:@39444.6]
  wire [31:0] _GEN_2109; // @[AxiLoadQueue.scala 268:32:@39438.4]
  wire [31:0] _GEN_2110; // @[AxiLoadQueue.scala 270:79:@39453.6]
  wire [31:0] _GEN_2111; // @[AxiLoadQueue.scala 268:32:@39447.4]
  wire [31:0] _GEN_2112; // @[AxiLoadQueue.scala 270:79:@39462.6]
  wire [31:0] _GEN_2113; // @[AxiLoadQueue.scala 268:32:@39456.4]
  wire [31:0] _GEN_2114; // @[AxiLoadQueue.scala 270:79:@39471.6]
  wire [31:0] _GEN_2115; // @[AxiLoadQueue.scala 268:32:@39465.4]
  wire [31:0] _GEN_2116; // @[AxiLoadQueue.scala 270:79:@39480.6]
  wire [31:0] _GEN_2117; // @[AxiLoadQueue.scala 268:32:@39474.4]
  wire [31:0] _GEN_2118; // @[AxiLoadQueue.scala 270:79:@39489.6]
  wire [31:0] _GEN_2119; // @[AxiLoadQueue.scala 268:32:@39483.4]
  wire [31:0] _GEN_2120; // @[AxiLoadQueue.scala 270:79:@39498.6]
  wire [31:0] _GEN_2121; // @[AxiLoadQueue.scala 268:32:@39492.4]
  wire [31:0] _GEN_2122; // @[AxiLoadQueue.scala 270:79:@39507.6]
  wire [31:0] _GEN_2123; // @[AxiLoadQueue.scala 268:32:@39501.4]
  wire [31:0] _GEN_2124; // @[AxiLoadQueue.scala 270:79:@39516.6]
  wire [31:0] _GEN_2125; // @[AxiLoadQueue.scala 268:32:@39510.4]
  wire [31:0] _GEN_2126; // @[AxiLoadQueue.scala 270:79:@39525.6]
  wire [31:0] _GEN_2127; // @[AxiLoadQueue.scala 268:32:@39519.4]
  wire  entriesPorts_0_0; // @[AxiLoadQueue.scala 288:69:@39529.4]
  wire  entriesPorts_0_1; // @[AxiLoadQueue.scala 288:69:@39531.4]
  wire  entriesPorts_0_2; // @[AxiLoadQueue.scala 288:69:@39533.4]
  wire  entriesPorts_0_3; // @[AxiLoadQueue.scala 288:69:@39535.4]
  wire  entriesPorts_0_4; // @[AxiLoadQueue.scala 288:69:@39537.4]
  wire  entriesPorts_0_5; // @[AxiLoadQueue.scala 288:69:@39539.4]
  wire  entriesPorts_0_6; // @[AxiLoadQueue.scala 288:69:@39541.4]
  wire  entriesPorts_0_7; // @[AxiLoadQueue.scala 288:69:@39543.4]
  wire  entriesPorts_0_8; // @[AxiLoadQueue.scala 288:69:@39545.4]
  wire  entriesPorts_0_9; // @[AxiLoadQueue.scala 288:69:@39547.4]
  wire  entriesPorts_0_10; // @[AxiLoadQueue.scala 288:69:@39549.4]
  wire  entriesPorts_0_11; // @[AxiLoadQueue.scala 288:69:@39551.4]
  wire  entriesPorts_0_12; // @[AxiLoadQueue.scala 288:69:@39553.4]
  wire  entriesPorts_0_13; // @[AxiLoadQueue.scala 288:69:@39555.4]
  wire  entriesPorts_0_14; // @[AxiLoadQueue.scala 288:69:@39557.4]
  wire  entriesPorts_0_15; // @[AxiLoadQueue.scala 288:69:@39559.4]
  wire  _T_94318; // @[AxiLoadQueue.scala 300:86:@39563.4]
  wire  _T_94319; // @[AxiLoadQueue.scala 300:83:@39564.4]
  wire  _T_94321; // @[AxiLoadQueue.scala 300:86:@39565.4]
  wire  _T_94322; // @[AxiLoadQueue.scala 300:83:@39566.4]
  wire  _T_94324; // @[AxiLoadQueue.scala 300:86:@39567.4]
  wire  _T_94325; // @[AxiLoadQueue.scala 300:83:@39568.4]
  wire  _T_94327; // @[AxiLoadQueue.scala 300:86:@39569.4]
  wire  _T_94328; // @[AxiLoadQueue.scala 300:83:@39570.4]
  wire  _T_94330; // @[AxiLoadQueue.scala 300:86:@39571.4]
  wire  _T_94331; // @[AxiLoadQueue.scala 300:83:@39572.4]
  wire  _T_94333; // @[AxiLoadQueue.scala 300:86:@39573.4]
  wire  _T_94334; // @[AxiLoadQueue.scala 300:83:@39574.4]
  wire  _T_94336; // @[AxiLoadQueue.scala 300:86:@39575.4]
  wire  _T_94337; // @[AxiLoadQueue.scala 300:83:@39576.4]
  wire  _T_94339; // @[AxiLoadQueue.scala 300:86:@39577.4]
  wire  _T_94340; // @[AxiLoadQueue.scala 300:83:@39578.4]
  wire  _T_94342; // @[AxiLoadQueue.scala 300:86:@39579.4]
  wire  _T_94343; // @[AxiLoadQueue.scala 300:83:@39580.4]
  wire  _T_94345; // @[AxiLoadQueue.scala 300:86:@39581.4]
  wire  _T_94346; // @[AxiLoadQueue.scala 300:83:@39582.4]
  wire  _T_94348; // @[AxiLoadQueue.scala 300:86:@39583.4]
  wire  _T_94349; // @[AxiLoadQueue.scala 300:83:@39584.4]
  wire  _T_94351; // @[AxiLoadQueue.scala 300:86:@39585.4]
  wire  _T_94352; // @[AxiLoadQueue.scala 300:83:@39586.4]
  wire  _T_94354; // @[AxiLoadQueue.scala 300:86:@39587.4]
  wire  _T_94355; // @[AxiLoadQueue.scala 300:83:@39588.4]
  wire  _T_94357; // @[AxiLoadQueue.scala 300:86:@39589.4]
  wire  _T_94358; // @[AxiLoadQueue.scala 300:83:@39590.4]
  wire  _T_94360; // @[AxiLoadQueue.scala 300:86:@39591.4]
  wire  _T_94361; // @[AxiLoadQueue.scala 300:83:@39592.4]
  wire  _T_94363; // @[AxiLoadQueue.scala 300:86:@39593.4]
  wire  _T_94364; // @[AxiLoadQueue.scala 300:83:@39594.4]
  wire [15:0] _T_94447; // @[Mux.scala 31:69:@39648.4]
  wire [15:0] _T_94448; // @[Mux.scala 31:69:@39649.4]
  wire [15:0] _T_94449; // @[Mux.scala 31:69:@39650.4]
  wire [15:0] _T_94450; // @[Mux.scala 31:69:@39651.4]
  wire [15:0] _T_94451; // @[Mux.scala 31:69:@39652.4]
  wire [15:0] _T_94452; // @[Mux.scala 31:69:@39653.4]
  wire [15:0] _T_94453; // @[Mux.scala 31:69:@39654.4]
  wire [15:0] _T_94454; // @[Mux.scala 31:69:@39655.4]
  wire [15:0] _T_94455; // @[Mux.scala 31:69:@39656.4]
  wire [15:0] _T_94456; // @[Mux.scala 31:69:@39657.4]
  wire [15:0] _T_94457; // @[Mux.scala 31:69:@39658.4]
  wire [15:0] _T_94458; // @[Mux.scala 31:69:@39659.4]
  wire [15:0] _T_94459; // @[Mux.scala 31:69:@39660.4]
  wire [15:0] _T_94460; // @[Mux.scala 31:69:@39661.4]
  wire [15:0] _T_94461; // @[Mux.scala 31:69:@39662.4]
  wire [15:0] _T_94462; // @[Mux.scala 31:69:@39663.4]
  wire  _T_94463; // @[OneHot.scala 66:30:@39664.4]
  wire  _T_94464; // @[OneHot.scala 66:30:@39665.4]
  wire  _T_94465; // @[OneHot.scala 66:30:@39666.4]
  wire  _T_94466; // @[OneHot.scala 66:30:@39667.4]
  wire  _T_94467; // @[OneHot.scala 66:30:@39668.4]
  wire  _T_94468; // @[OneHot.scala 66:30:@39669.4]
  wire  _T_94469; // @[OneHot.scala 66:30:@39670.4]
  wire  _T_94470; // @[OneHot.scala 66:30:@39671.4]
  wire  _T_94471; // @[OneHot.scala 66:30:@39672.4]
  wire  _T_94472; // @[OneHot.scala 66:30:@39673.4]
  wire  _T_94473; // @[OneHot.scala 66:30:@39674.4]
  wire  _T_94474; // @[OneHot.scala 66:30:@39675.4]
  wire  _T_94475; // @[OneHot.scala 66:30:@39676.4]
  wire  _T_94476; // @[OneHot.scala 66:30:@39677.4]
  wire  _T_94477; // @[OneHot.scala 66:30:@39678.4]
  wire  _T_94478; // @[OneHot.scala 66:30:@39679.4]
  wire [15:0] _T_94519; // @[Mux.scala 31:69:@39697.4]
  wire [15:0] _T_94520; // @[Mux.scala 31:69:@39698.4]
  wire [15:0] _T_94521; // @[Mux.scala 31:69:@39699.4]
  wire [15:0] _T_94522; // @[Mux.scala 31:69:@39700.4]
  wire [15:0] _T_94523; // @[Mux.scala 31:69:@39701.4]
  wire [15:0] _T_94524; // @[Mux.scala 31:69:@39702.4]
  wire [15:0] _T_94525; // @[Mux.scala 31:69:@39703.4]
  wire [15:0] _T_94526; // @[Mux.scala 31:69:@39704.4]
  wire [15:0] _T_94527; // @[Mux.scala 31:69:@39705.4]
  wire [15:0] _T_94528; // @[Mux.scala 31:69:@39706.4]
  wire [15:0] _T_94529; // @[Mux.scala 31:69:@39707.4]
  wire [15:0] _T_94530; // @[Mux.scala 31:69:@39708.4]
  wire [15:0] _T_94531; // @[Mux.scala 31:69:@39709.4]
  wire [15:0] _T_94532; // @[Mux.scala 31:69:@39710.4]
  wire [15:0] _T_94533; // @[Mux.scala 31:69:@39711.4]
  wire [15:0] _T_94534; // @[Mux.scala 31:69:@39712.4]
  wire  _T_94535; // @[OneHot.scala 66:30:@39713.4]
  wire  _T_94536; // @[OneHot.scala 66:30:@39714.4]
  wire  _T_94537; // @[OneHot.scala 66:30:@39715.4]
  wire  _T_94538; // @[OneHot.scala 66:30:@39716.4]
  wire  _T_94539; // @[OneHot.scala 66:30:@39717.4]
  wire  _T_94540; // @[OneHot.scala 66:30:@39718.4]
  wire  _T_94541; // @[OneHot.scala 66:30:@39719.4]
  wire  _T_94542; // @[OneHot.scala 66:30:@39720.4]
  wire  _T_94543; // @[OneHot.scala 66:30:@39721.4]
  wire  _T_94544; // @[OneHot.scala 66:30:@39722.4]
  wire  _T_94545; // @[OneHot.scala 66:30:@39723.4]
  wire  _T_94546; // @[OneHot.scala 66:30:@39724.4]
  wire  _T_94547; // @[OneHot.scala 66:30:@39725.4]
  wire  _T_94548; // @[OneHot.scala 66:30:@39726.4]
  wire  _T_94549; // @[OneHot.scala 66:30:@39727.4]
  wire  _T_94550; // @[OneHot.scala 66:30:@39728.4]
  wire [15:0] _T_94591; // @[Mux.scala 31:69:@39746.4]
  wire [15:0] _T_94592; // @[Mux.scala 31:69:@39747.4]
  wire [15:0] _T_94593; // @[Mux.scala 31:69:@39748.4]
  wire [15:0] _T_94594; // @[Mux.scala 31:69:@39749.4]
  wire [15:0] _T_94595; // @[Mux.scala 31:69:@39750.4]
  wire [15:0] _T_94596; // @[Mux.scala 31:69:@39751.4]
  wire [15:0] _T_94597; // @[Mux.scala 31:69:@39752.4]
  wire [15:0] _T_94598; // @[Mux.scala 31:69:@39753.4]
  wire [15:0] _T_94599; // @[Mux.scala 31:69:@39754.4]
  wire [15:0] _T_94600; // @[Mux.scala 31:69:@39755.4]
  wire [15:0] _T_94601; // @[Mux.scala 31:69:@39756.4]
  wire [15:0] _T_94602; // @[Mux.scala 31:69:@39757.4]
  wire [15:0] _T_94603; // @[Mux.scala 31:69:@39758.4]
  wire [15:0] _T_94604; // @[Mux.scala 31:69:@39759.4]
  wire [15:0] _T_94605; // @[Mux.scala 31:69:@39760.4]
  wire [15:0] _T_94606; // @[Mux.scala 31:69:@39761.4]
  wire  _T_94607; // @[OneHot.scala 66:30:@39762.4]
  wire  _T_94608; // @[OneHot.scala 66:30:@39763.4]
  wire  _T_94609; // @[OneHot.scala 66:30:@39764.4]
  wire  _T_94610; // @[OneHot.scala 66:30:@39765.4]
  wire  _T_94611; // @[OneHot.scala 66:30:@39766.4]
  wire  _T_94612; // @[OneHot.scala 66:30:@39767.4]
  wire  _T_94613; // @[OneHot.scala 66:30:@39768.4]
  wire  _T_94614; // @[OneHot.scala 66:30:@39769.4]
  wire  _T_94615; // @[OneHot.scala 66:30:@39770.4]
  wire  _T_94616; // @[OneHot.scala 66:30:@39771.4]
  wire  _T_94617; // @[OneHot.scala 66:30:@39772.4]
  wire  _T_94618; // @[OneHot.scala 66:30:@39773.4]
  wire  _T_94619; // @[OneHot.scala 66:30:@39774.4]
  wire  _T_94620; // @[OneHot.scala 66:30:@39775.4]
  wire  _T_94621; // @[OneHot.scala 66:30:@39776.4]
  wire  _T_94622; // @[OneHot.scala 66:30:@39777.4]
  wire [15:0] _T_94663; // @[Mux.scala 31:69:@39795.4]
  wire [15:0] _T_94664; // @[Mux.scala 31:69:@39796.4]
  wire [15:0] _T_94665; // @[Mux.scala 31:69:@39797.4]
  wire [15:0] _T_94666; // @[Mux.scala 31:69:@39798.4]
  wire [15:0] _T_94667; // @[Mux.scala 31:69:@39799.4]
  wire [15:0] _T_94668; // @[Mux.scala 31:69:@39800.4]
  wire [15:0] _T_94669; // @[Mux.scala 31:69:@39801.4]
  wire [15:0] _T_94670; // @[Mux.scala 31:69:@39802.4]
  wire [15:0] _T_94671; // @[Mux.scala 31:69:@39803.4]
  wire [15:0] _T_94672; // @[Mux.scala 31:69:@39804.4]
  wire [15:0] _T_94673; // @[Mux.scala 31:69:@39805.4]
  wire [15:0] _T_94674; // @[Mux.scala 31:69:@39806.4]
  wire [15:0] _T_94675; // @[Mux.scala 31:69:@39807.4]
  wire [15:0] _T_94676; // @[Mux.scala 31:69:@39808.4]
  wire [15:0] _T_94677; // @[Mux.scala 31:69:@39809.4]
  wire [15:0] _T_94678; // @[Mux.scala 31:69:@39810.4]
  wire  _T_94679; // @[OneHot.scala 66:30:@39811.4]
  wire  _T_94680; // @[OneHot.scala 66:30:@39812.4]
  wire  _T_94681; // @[OneHot.scala 66:30:@39813.4]
  wire  _T_94682; // @[OneHot.scala 66:30:@39814.4]
  wire  _T_94683; // @[OneHot.scala 66:30:@39815.4]
  wire  _T_94684; // @[OneHot.scala 66:30:@39816.4]
  wire  _T_94685; // @[OneHot.scala 66:30:@39817.4]
  wire  _T_94686; // @[OneHot.scala 66:30:@39818.4]
  wire  _T_94687; // @[OneHot.scala 66:30:@39819.4]
  wire  _T_94688; // @[OneHot.scala 66:30:@39820.4]
  wire  _T_94689; // @[OneHot.scala 66:30:@39821.4]
  wire  _T_94690; // @[OneHot.scala 66:30:@39822.4]
  wire  _T_94691; // @[OneHot.scala 66:30:@39823.4]
  wire  _T_94692; // @[OneHot.scala 66:30:@39824.4]
  wire  _T_94693; // @[OneHot.scala 66:30:@39825.4]
  wire  _T_94694; // @[OneHot.scala 66:30:@39826.4]
  wire [15:0] _T_94735; // @[Mux.scala 31:69:@39844.4]
  wire [15:0] _T_94736; // @[Mux.scala 31:69:@39845.4]
  wire [15:0] _T_94737; // @[Mux.scala 31:69:@39846.4]
  wire [15:0] _T_94738; // @[Mux.scala 31:69:@39847.4]
  wire [15:0] _T_94739; // @[Mux.scala 31:69:@39848.4]
  wire [15:0] _T_94740; // @[Mux.scala 31:69:@39849.4]
  wire [15:0] _T_94741; // @[Mux.scala 31:69:@39850.4]
  wire [15:0] _T_94742; // @[Mux.scala 31:69:@39851.4]
  wire [15:0] _T_94743; // @[Mux.scala 31:69:@39852.4]
  wire [15:0] _T_94744; // @[Mux.scala 31:69:@39853.4]
  wire [15:0] _T_94745; // @[Mux.scala 31:69:@39854.4]
  wire [15:0] _T_94746; // @[Mux.scala 31:69:@39855.4]
  wire [15:0] _T_94747; // @[Mux.scala 31:69:@39856.4]
  wire [15:0] _T_94748; // @[Mux.scala 31:69:@39857.4]
  wire [15:0] _T_94749; // @[Mux.scala 31:69:@39858.4]
  wire [15:0] _T_94750; // @[Mux.scala 31:69:@39859.4]
  wire  _T_94751; // @[OneHot.scala 66:30:@39860.4]
  wire  _T_94752; // @[OneHot.scala 66:30:@39861.4]
  wire  _T_94753; // @[OneHot.scala 66:30:@39862.4]
  wire  _T_94754; // @[OneHot.scala 66:30:@39863.4]
  wire  _T_94755; // @[OneHot.scala 66:30:@39864.4]
  wire  _T_94756; // @[OneHot.scala 66:30:@39865.4]
  wire  _T_94757; // @[OneHot.scala 66:30:@39866.4]
  wire  _T_94758; // @[OneHot.scala 66:30:@39867.4]
  wire  _T_94759; // @[OneHot.scala 66:30:@39868.4]
  wire  _T_94760; // @[OneHot.scala 66:30:@39869.4]
  wire  _T_94761; // @[OneHot.scala 66:30:@39870.4]
  wire  _T_94762; // @[OneHot.scala 66:30:@39871.4]
  wire  _T_94763; // @[OneHot.scala 66:30:@39872.4]
  wire  _T_94764; // @[OneHot.scala 66:30:@39873.4]
  wire  _T_94765; // @[OneHot.scala 66:30:@39874.4]
  wire  _T_94766; // @[OneHot.scala 66:30:@39875.4]
  wire [15:0] _T_94807; // @[Mux.scala 31:69:@39893.4]
  wire [15:0] _T_94808; // @[Mux.scala 31:69:@39894.4]
  wire [15:0] _T_94809; // @[Mux.scala 31:69:@39895.4]
  wire [15:0] _T_94810; // @[Mux.scala 31:69:@39896.4]
  wire [15:0] _T_94811; // @[Mux.scala 31:69:@39897.4]
  wire [15:0] _T_94812; // @[Mux.scala 31:69:@39898.4]
  wire [15:0] _T_94813; // @[Mux.scala 31:69:@39899.4]
  wire [15:0] _T_94814; // @[Mux.scala 31:69:@39900.4]
  wire [15:0] _T_94815; // @[Mux.scala 31:69:@39901.4]
  wire [15:0] _T_94816; // @[Mux.scala 31:69:@39902.4]
  wire [15:0] _T_94817; // @[Mux.scala 31:69:@39903.4]
  wire [15:0] _T_94818; // @[Mux.scala 31:69:@39904.4]
  wire [15:0] _T_94819; // @[Mux.scala 31:69:@39905.4]
  wire [15:0] _T_94820; // @[Mux.scala 31:69:@39906.4]
  wire [15:0] _T_94821; // @[Mux.scala 31:69:@39907.4]
  wire [15:0] _T_94822; // @[Mux.scala 31:69:@39908.4]
  wire  _T_94823; // @[OneHot.scala 66:30:@39909.4]
  wire  _T_94824; // @[OneHot.scala 66:30:@39910.4]
  wire  _T_94825; // @[OneHot.scala 66:30:@39911.4]
  wire  _T_94826; // @[OneHot.scala 66:30:@39912.4]
  wire  _T_94827; // @[OneHot.scala 66:30:@39913.4]
  wire  _T_94828; // @[OneHot.scala 66:30:@39914.4]
  wire  _T_94829; // @[OneHot.scala 66:30:@39915.4]
  wire  _T_94830; // @[OneHot.scala 66:30:@39916.4]
  wire  _T_94831; // @[OneHot.scala 66:30:@39917.4]
  wire  _T_94832; // @[OneHot.scala 66:30:@39918.4]
  wire  _T_94833; // @[OneHot.scala 66:30:@39919.4]
  wire  _T_94834; // @[OneHot.scala 66:30:@39920.4]
  wire  _T_94835; // @[OneHot.scala 66:30:@39921.4]
  wire  _T_94836; // @[OneHot.scala 66:30:@39922.4]
  wire  _T_94837; // @[OneHot.scala 66:30:@39923.4]
  wire  _T_94838; // @[OneHot.scala 66:30:@39924.4]
  wire [15:0] _T_94879; // @[Mux.scala 31:69:@39942.4]
  wire [15:0] _T_94880; // @[Mux.scala 31:69:@39943.4]
  wire [15:0] _T_94881; // @[Mux.scala 31:69:@39944.4]
  wire [15:0] _T_94882; // @[Mux.scala 31:69:@39945.4]
  wire [15:0] _T_94883; // @[Mux.scala 31:69:@39946.4]
  wire [15:0] _T_94884; // @[Mux.scala 31:69:@39947.4]
  wire [15:0] _T_94885; // @[Mux.scala 31:69:@39948.4]
  wire [15:0] _T_94886; // @[Mux.scala 31:69:@39949.4]
  wire [15:0] _T_94887; // @[Mux.scala 31:69:@39950.4]
  wire [15:0] _T_94888; // @[Mux.scala 31:69:@39951.4]
  wire [15:0] _T_94889; // @[Mux.scala 31:69:@39952.4]
  wire [15:0] _T_94890; // @[Mux.scala 31:69:@39953.4]
  wire [15:0] _T_94891; // @[Mux.scala 31:69:@39954.4]
  wire [15:0] _T_94892; // @[Mux.scala 31:69:@39955.4]
  wire [15:0] _T_94893; // @[Mux.scala 31:69:@39956.4]
  wire [15:0] _T_94894; // @[Mux.scala 31:69:@39957.4]
  wire  _T_94895; // @[OneHot.scala 66:30:@39958.4]
  wire  _T_94896; // @[OneHot.scala 66:30:@39959.4]
  wire  _T_94897; // @[OneHot.scala 66:30:@39960.4]
  wire  _T_94898; // @[OneHot.scala 66:30:@39961.4]
  wire  _T_94899; // @[OneHot.scala 66:30:@39962.4]
  wire  _T_94900; // @[OneHot.scala 66:30:@39963.4]
  wire  _T_94901; // @[OneHot.scala 66:30:@39964.4]
  wire  _T_94902; // @[OneHot.scala 66:30:@39965.4]
  wire  _T_94903; // @[OneHot.scala 66:30:@39966.4]
  wire  _T_94904; // @[OneHot.scala 66:30:@39967.4]
  wire  _T_94905; // @[OneHot.scala 66:30:@39968.4]
  wire  _T_94906; // @[OneHot.scala 66:30:@39969.4]
  wire  _T_94907; // @[OneHot.scala 66:30:@39970.4]
  wire  _T_94908; // @[OneHot.scala 66:30:@39971.4]
  wire  _T_94909; // @[OneHot.scala 66:30:@39972.4]
  wire  _T_94910; // @[OneHot.scala 66:30:@39973.4]
  wire [15:0] _T_94951; // @[Mux.scala 31:69:@39991.4]
  wire [15:0] _T_94952; // @[Mux.scala 31:69:@39992.4]
  wire [15:0] _T_94953; // @[Mux.scala 31:69:@39993.4]
  wire [15:0] _T_94954; // @[Mux.scala 31:69:@39994.4]
  wire [15:0] _T_94955; // @[Mux.scala 31:69:@39995.4]
  wire [15:0] _T_94956; // @[Mux.scala 31:69:@39996.4]
  wire [15:0] _T_94957; // @[Mux.scala 31:69:@39997.4]
  wire [15:0] _T_94958; // @[Mux.scala 31:69:@39998.4]
  wire [15:0] _T_94959; // @[Mux.scala 31:69:@39999.4]
  wire [15:0] _T_94960; // @[Mux.scala 31:69:@40000.4]
  wire [15:0] _T_94961; // @[Mux.scala 31:69:@40001.4]
  wire [15:0] _T_94962; // @[Mux.scala 31:69:@40002.4]
  wire [15:0] _T_94963; // @[Mux.scala 31:69:@40003.4]
  wire [15:0] _T_94964; // @[Mux.scala 31:69:@40004.4]
  wire [15:0] _T_94965; // @[Mux.scala 31:69:@40005.4]
  wire [15:0] _T_94966; // @[Mux.scala 31:69:@40006.4]
  wire  _T_94967; // @[OneHot.scala 66:30:@40007.4]
  wire  _T_94968; // @[OneHot.scala 66:30:@40008.4]
  wire  _T_94969; // @[OneHot.scala 66:30:@40009.4]
  wire  _T_94970; // @[OneHot.scala 66:30:@40010.4]
  wire  _T_94971; // @[OneHot.scala 66:30:@40011.4]
  wire  _T_94972; // @[OneHot.scala 66:30:@40012.4]
  wire  _T_94973; // @[OneHot.scala 66:30:@40013.4]
  wire  _T_94974; // @[OneHot.scala 66:30:@40014.4]
  wire  _T_94975; // @[OneHot.scala 66:30:@40015.4]
  wire  _T_94976; // @[OneHot.scala 66:30:@40016.4]
  wire  _T_94977; // @[OneHot.scala 66:30:@40017.4]
  wire  _T_94978; // @[OneHot.scala 66:30:@40018.4]
  wire  _T_94979; // @[OneHot.scala 66:30:@40019.4]
  wire  _T_94980; // @[OneHot.scala 66:30:@40020.4]
  wire  _T_94981; // @[OneHot.scala 66:30:@40021.4]
  wire  _T_94982; // @[OneHot.scala 66:30:@40022.4]
  wire [15:0] _T_95023; // @[Mux.scala 31:69:@40040.4]
  wire [15:0] _T_95024; // @[Mux.scala 31:69:@40041.4]
  wire [15:0] _T_95025; // @[Mux.scala 31:69:@40042.4]
  wire [15:0] _T_95026; // @[Mux.scala 31:69:@40043.4]
  wire [15:0] _T_95027; // @[Mux.scala 31:69:@40044.4]
  wire [15:0] _T_95028; // @[Mux.scala 31:69:@40045.4]
  wire [15:0] _T_95029; // @[Mux.scala 31:69:@40046.4]
  wire [15:0] _T_95030; // @[Mux.scala 31:69:@40047.4]
  wire [15:0] _T_95031; // @[Mux.scala 31:69:@40048.4]
  wire [15:0] _T_95032; // @[Mux.scala 31:69:@40049.4]
  wire [15:0] _T_95033; // @[Mux.scala 31:69:@40050.4]
  wire [15:0] _T_95034; // @[Mux.scala 31:69:@40051.4]
  wire [15:0] _T_95035; // @[Mux.scala 31:69:@40052.4]
  wire [15:0] _T_95036; // @[Mux.scala 31:69:@40053.4]
  wire [15:0] _T_95037; // @[Mux.scala 31:69:@40054.4]
  wire [15:0] _T_95038; // @[Mux.scala 31:69:@40055.4]
  wire  _T_95039; // @[OneHot.scala 66:30:@40056.4]
  wire  _T_95040; // @[OneHot.scala 66:30:@40057.4]
  wire  _T_95041; // @[OneHot.scala 66:30:@40058.4]
  wire  _T_95042; // @[OneHot.scala 66:30:@40059.4]
  wire  _T_95043; // @[OneHot.scala 66:30:@40060.4]
  wire  _T_95044; // @[OneHot.scala 66:30:@40061.4]
  wire  _T_95045; // @[OneHot.scala 66:30:@40062.4]
  wire  _T_95046; // @[OneHot.scala 66:30:@40063.4]
  wire  _T_95047; // @[OneHot.scala 66:30:@40064.4]
  wire  _T_95048; // @[OneHot.scala 66:30:@40065.4]
  wire  _T_95049; // @[OneHot.scala 66:30:@40066.4]
  wire  _T_95050; // @[OneHot.scala 66:30:@40067.4]
  wire  _T_95051; // @[OneHot.scala 66:30:@40068.4]
  wire  _T_95052; // @[OneHot.scala 66:30:@40069.4]
  wire  _T_95053; // @[OneHot.scala 66:30:@40070.4]
  wire  _T_95054; // @[OneHot.scala 66:30:@40071.4]
  wire [15:0] _T_95095; // @[Mux.scala 31:69:@40089.4]
  wire [15:0] _T_95096; // @[Mux.scala 31:69:@40090.4]
  wire [15:0] _T_95097; // @[Mux.scala 31:69:@40091.4]
  wire [15:0] _T_95098; // @[Mux.scala 31:69:@40092.4]
  wire [15:0] _T_95099; // @[Mux.scala 31:69:@40093.4]
  wire [15:0] _T_95100; // @[Mux.scala 31:69:@40094.4]
  wire [15:0] _T_95101; // @[Mux.scala 31:69:@40095.4]
  wire [15:0] _T_95102; // @[Mux.scala 31:69:@40096.4]
  wire [15:0] _T_95103; // @[Mux.scala 31:69:@40097.4]
  wire [15:0] _T_95104; // @[Mux.scala 31:69:@40098.4]
  wire [15:0] _T_95105; // @[Mux.scala 31:69:@40099.4]
  wire [15:0] _T_95106; // @[Mux.scala 31:69:@40100.4]
  wire [15:0] _T_95107; // @[Mux.scala 31:69:@40101.4]
  wire [15:0] _T_95108; // @[Mux.scala 31:69:@40102.4]
  wire [15:0] _T_95109; // @[Mux.scala 31:69:@40103.4]
  wire [15:0] _T_95110; // @[Mux.scala 31:69:@40104.4]
  wire  _T_95111; // @[OneHot.scala 66:30:@40105.4]
  wire  _T_95112; // @[OneHot.scala 66:30:@40106.4]
  wire  _T_95113; // @[OneHot.scala 66:30:@40107.4]
  wire  _T_95114; // @[OneHot.scala 66:30:@40108.4]
  wire  _T_95115; // @[OneHot.scala 66:30:@40109.4]
  wire  _T_95116; // @[OneHot.scala 66:30:@40110.4]
  wire  _T_95117; // @[OneHot.scala 66:30:@40111.4]
  wire  _T_95118; // @[OneHot.scala 66:30:@40112.4]
  wire  _T_95119; // @[OneHot.scala 66:30:@40113.4]
  wire  _T_95120; // @[OneHot.scala 66:30:@40114.4]
  wire  _T_95121; // @[OneHot.scala 66:30:@40115.4]
  wire  _T_95122; // @[OneHot.scala 66:30:@40116.4]
  wire  _T_95123; // @[OneHot.scala 66:30:@40117.4]
  wire  _T_95124; // @[OneHot.scala 66:30:@40118.4]
  wire  _T_95125; // @[OneHot.scala 66:30:@40119.4]
  wire  _T_95126; // @[OneHot.scala 66:30:@40120.4]
  wire [15:0] _T_95167; // @[Mux.scala 31:69:@40138.4]
  wire [15:0] _T_95168; // @[Mux.scala 31:69:@40139.4]
  wire [15:0] _T_95169; // @[Mux.scala 31:69:@40140.4]
  wire [15:0] _T_95170; // @[Mux.scala 31:69:@40141.4]
  wire [15:0] _T_95171; // @[Mux.scala 31:69:@40142.4]
  wire [15:0] _T_95172; // @[Mux.scala 31:69:@40143.4]
  wire [15:0] _T_95173; // @[Mux.scala 31:69:@40144.4]
  wire [15:0] _T_95174; // @[Mux.scala 31:69:@40145.4]
  wire [15:0] _T_95175; // @[Mux.scala 31:69:@40146.4]
  wire [15:0] _T_95176; // @[Mux.scala 31:69:@40147.4]
  wire [15:0] _T_95177; // @[Mux.scala 31:69:@40148.4]
  wire [15:0] _T_95178; // @[Mux.scala 31:69:@40149.4]
  wire [15:0] _T_95179; // @[Mux.scala 31:69:@40150.4]
  wire [15:0] _T_95180; // @[Mux.scala 31:69:@40151.4]
  wire [15:0] _T_95181; // @[Mux.scala 31:69:@40152.4]
  wire [15:0] _T_95182; // @[Mux.scala 31:69:@40153.4]
  wire  _T_95183; // @[OneHot.scala 66:30:@40154.4]
  wire  _T_95184; // @[OneHot.scala 66:30:@40155.4]
  wire  _T_95185; // @[OneHot.scala 66:30:@40156.4]
  wire  _T_95186; // @[OneHot.scala 66:30:@40157.4]
  wire  _T_95187; // @[OneHot.scala 66:30:@40158.4]
  wire  _T_95188; // @[OneHot.scala 66:30:@40159.4]
  wire  _T_95189; // @[OneHot.scala 66:30:@40160.4]
  wire  _T_95190; // @[OneHot.scala 66:30:@40161.4]
  wire  _T_95191; // @[OneHot.scala 66:30:@40162.4]
  wire  _T_95192; // @[OneHot.scala 66:30:@40163.4]
  wire  _T_95193; // @[OneHot.scala 66:30:@40164.4]
  wire  _T_95194; // @[OneHot.scala 66:30:@40165.4]
  wire  _T_95195; // @[OneHot.scala 66:30:@40166.4]
  wire  _T_95196; // @[OneHot.scala 66:30:@40167.4]
  wire  _T_95197; // @[OneHot.scala 66:30:@40168.4]
  wire  _T_95198; // @[OneHot.scala 66:30:@40169.4]
  wire [15:0] _T_95239; // @[Mux.scala 31:69:@40187.4]
  wire [15:0] _T_95240; // @[Mux.scala 31:69:@40188.4]
  wire [15:0] _T_95241; // @[Mux.scala 31:69:@40189.4]
  wire [15:0] _T_95242; // @[Mux.scala 31:69:@40190.4]
  wire [15:0] _T_95243; // @[Mux.scala 31:69:@40191.4]
  wire [15:0] _T_95244; // @[Mux.scala 31:69:@40192.4]
  wire [15:0] _T_95245; // @[Mux.scala 31:69:@40193.4]
  wire [15:0] _T_95246; // @[Mux.scala 31:69:@40194.4]
  wire [15:0] _T_95247; // @[Mux.scala 31:69:@40195.4]
  wire [15:0] _T_95248; // @[Mux.scala 31:69:@40196.4]
  wire [15:0] _T_95249; // @[Mux.scala 31:69:@40197.4]
  wire [15:0] _T_95250; // @[Mux.scala 31:69:@40198.4]
  wire [15:0] _T_95251; // @[Mux.scala 31:69:@40199.4]
  wire [15:0] _T_95252; // @[Mux.scala 31:69:@40200.4]
  wire [15:0] _T_95253; // @[Mux.scala 31:69:@40201.4]
  wire [15:0] _T_95254; // @[Mux.scala 31:69:@40202.4]
  wire  _T_95255; // @[OneHot.scala 66:30:@40203.4]
  wire  _T_95256; // @[OneHot.scala 66:30:@40204.4]
  wire  _T_95257; // @[OneHot.scala 66:30:@40205.4]
  wire  _T_95258; // @[OneHot.scala 66:30:@40206.4]
  wire  _T_95259; // @[OneHot.scala 66:30:@40207.4]
  wire  _T_95260; // @[OneHot.scala 66:30:@40208.4]
  wire  _T_95261; // @[OneHot.scala 66:30:@40209.4]
  wire  _T_95262; // @[OneHot.scala 66:30:@40210.4]
  wire  _T_95263; // @[OneHot.scala 66:30:@40211.4]
  wire  _T_95264; // @[OneHot.scala 66:30:@40212.4]
  wire  _T_95265; // @[OneHot.scala 66:30:@40213.4]
  wire  _T_95266; // @[OneHot.scala 66:30:@40214.4]
  wire  _T_95267; // @[OneHot.scala 66:30:@40215.4]
  wire  _T_95268; // @[OneHot.scala 66:30:@40216.4]
  wire  _T_95269; // @[OneHot.scala 66:30:@40217.4]
  wire  _T_95270; // @[OneHot.scala 66:30:@40218.4]
  wire [15:0] _T_95311; // @[Mux.scala 31:69:@40236.4]
  wire [15:0] _T_95312; // @[Mux.scala 31:69:@40237.4]
  wire [15:0] _T_95313; // @[Mux.scala 31:69:@40238.4]
  wire [15:0] _T_95314; // @[Mux.scala 31:69:@40239.4]
  wire [15:0] _T_95315; // @[Mux.scala 31:69:@40240.4]
  wire [15:0] _T_95316; // @[Mux.scala 31:69:@40241.4]
  wire [15:0] _T_95317; // @[Mux.scala 31:69:@40242.4]
  wire [15:0] _T_95318; // @[Mux.scala 31:69:@40243.4]
  wire [15:0] _T_95319; // @[Mux.scala 31:69:@40244.4]
  wire [15:0] _T_95320; // @[Mux.scala 31:69:@40245.4]
  wire [15:0] _T_95321; // @[Mux.scala 31:69:@40246.4]
  wire [15:0] _T_95322; // @[Mux.scala 31:69:@40247.4]
  wire [15:0] _T_95323; // @[Mux.scala 31:69:@40248.4]
  wire [15:0] _T_95324; // @[Mux.scala 31:69:@40249.4]
  wire [15:0] _T_95325; // @[Mux.scala 31:69:@40250.4]
  wire [15:0] _T_95326; // @[Mux.scala 31:69:@40251.4]
  wire  _T_95327; // @[OneHot.scala 66:30:@40252.4]
  wire  _T_95328; // @[OneHot.scala 66:30:@40253.4]
  wire  _T_95329; // @[OneHot.scala 66:30:@40254.4]
  wire  _T_95330; // @[OneHot.scala 66:30:@40255.4]
  wire  _T_95331; // @[OneHot.scala 66:30:@40256.4]
  wire  _T_95332; // @[OneHot.scala 66:30:@40257.4]
  wire  _T_95333; // @[OneHot.scala 66:30:@40258.4]
  wire  _T_95334; // @[OneHot.scala 66:30:@40259.4]
  wire  _T_95335; // @[OneHot.scala 66:30:@40260.4]
  wire  _T_95336; // @[OneHot.scala 66:30:@40261.4]
  wire  _T_95337; // @[OneHot.scala 66:30:@40262.4]
  wire  _T_95338; // @[OneHot.scala 66:30:@40263.4]
  wire  _T_95339; // @[OneHot.scala 66:30:@40264.4]
  wire  _T_95340; // @[OneHot.scala 66:30:@40265.4]
  wire  _T_95341; // @[OneHot.scala 66:30:@40266.4]
  wire  _T_95342; // @[OneHot.scala 66:30:@40267.4]
  wire [15:0] _T_95383; // @[Mux.scala 31:69:@40285.4]
  wire [15:0] _T_95384; // @[Mux.scala 31:69:@40286.4]
  wire [15:0] _T_95385; // @[Mux.scala 31:69:@40287.4]
  wire [15:0] _T_95386; // @[Mux.scala 31:69:@40288.4]
  wire [15:0] _T_95387; // @[Mux.scala 31:69:@40289.4]
  wire [15:0] _T_95388; // @[Mux.scala 31:69:@40290.4]
  wire [15:0] _T_95389; // @[Mux.scala 31:69:@40291.4]
  wire [15:0] _T_95390; // @[Mux.scala 31:69:@40292.4]
  wire [15:0] _T_95391; // @[Mux.scala 31:69:@40293.4]
  wire [15:0] _T_95392; // @[Mux.scala 31:69:@40294.4]
  wire [15:0] _T_95393; // @[Mux.scala 31:69:@40295.4]
  wire [15:0] _T_95394; // @[Mux.scala 31:69:@40296.4]
  wire [15:0] _T_95395; // @[Mux.scala 31:69:@40297.4]
  wire [15:0] _T_95396; // @[Mux.scala 31:69:@40298.4]
  wire [15:0] _T_95397; // @[Mux.scala 31:69:@40299.4]
  wire [15:0] _T_95398; // @[Mux.scala 31:69:@40300.4]
  wire  _T_95399; // @[OneHot.scala 66:30:@40301.4]
  wire  _T_95400; // @[OneHot.scala 66:30:@40302.4]
  wire  _T_95401; // @[OneHot.scala 66:30:@40303.4]
  wire  _T_95402; // @[OneHot.scala 66:30:@40304.4]
  wire  _T_95403; // @[OneHot.scala 66:30:@40305.4]
  wire  _T_95404; // @[OneHot.scala 66:30:@40306.4]
  wire  _T_95405; // @[OneHot.scala 66:30:@40307.4]
  wire  _T_95406; // @[OneHot.scala 66:30:@40308.4]
  wire  _T_95407; // @[OneHot.scala 66:30:@40309.4]
  wire  _T_95408; // @[OneHot.scala 66:30:@40310.4]
  wire  _T_95409; // @[OneHot.scala 66:30:@40311.4]
  wire  _T_95410; // @[OneHot.scala 66:30:@40312.4]
  wire  _T_95411; // @[OneHot.scala 66:30:@40313.4]
  wire  _T_95412; // @[OneHot.scala 66:30:@40314.4]
  wire  _T_95413; // @[OneHot.scala 66:30:@40315.4]
  wire  _T_95414; // @[OneHot.scala 66:30:@40316.4]
  wire [15:0] _T_95455; // @[Mux.scala 31:69:@40334.4]
  wire [15:0] _T_95456; // @[Mux.scala 31:69:@40335.4]
  wire [15:0] _T_95457; // @[Mux.scala 31:69:@40336.4]
  wire [15:0] _T_95458; // @[Mux.scala 31:69:@40337.4]
  wire [15:0] _T_95459; // @[Mux.scala 31:69:@40338.4]
  wire [15:0] _T_95460; // @[Mux.scala 31:69:@40339.4]
  wire [15:0] _T_95461; // @[Mux.scala 31:69:@40340.4]
  wire [15:0] _T_95462; // @[Mux.scala 31:69:@40341.4]
  wire [15:0] _T_95463; // @[Mux.scala 31:69:@40342.4]
  wire [15:0] _T_95464; // @[Mux.scala 31:69:@40343.4]
  wire [15:0] _T_95465; // @[Mux.scala 31:69:@40344.4]
  wire [15:0] _T_95466; // @[Mux.scala 31:69:@40345.4]
  wire [15:0] _T_95467; // @[Mux.scala 31:69:@40346.4]
  wire [15:0] _T_95468; // @[Mux.scala 31:69:@40347.4]
  wire [15:0] _T_95469; // @[Mux.scala 31:69:@40348.4]
  wire [15:0] _T_95470; // @[Mux.scala 31:69:@40349.4]
  wire  _T_95471; // @[OneHot.scala 66:30:@40350.4]
  wire  _T_95472; // @[OneHot.scala 66:30:@40351.4]
  wire  _T_95473; // @[OneHot.scala 66:30:@40352.4]
  wire  _T_95474; // @[OneHot.scala 66:30:@40353.4]
  wire  _T_95475; // @[OneHot.scala 66:30:@40354.4]
  wire  _T_95476; // @[OneHot.scala 66:30:@40355.4]
  wire  _T_95477; // @[OneHot.scala 66:30:@40356.4]
  wire  _T_95478; // @[OneHot.scala 66:30:@40357.4]
  wire  _T_95479; // @[OneHot.scala 66:30:@40358.4]
  wire  _T_95480; // @[OneHot.scala 66:30:@40359.4]
  wire  _T_95481; // @[OneHot.scala 66:30:@40360.4]
  wire  _T_95482; // @[OneHot.scala 66:30:@40361.4]
  wire  _T_95483; // @[OneHot.scala 66:30:@40362.4]
  wire  _T_95484; // @[OneHot.scala 66:30:@40363.4]
  wire  _T_95485; // @[OneHot.scala 66:30:@40364.4]
  wire  _T_95486; // @[OneHot.scala 66:30:@40365.4]
  wire [15:0] _T_95527; // @[Mux.scala 31:69:@40383.4]
  wire [15:0] _T_95528; // @[Mux.scala 31:69:@40384.4]
  wire [15:0] _T_95529; // @[Mux.scala 31:69:@40385.4]
  wire [15:0] _T_95530; // @[Mux.scala 31:69:@40386.4]
  wire [15:0] _T_95531; // @[Mux.scala 31:69:@40387.4]
  wire [15:0] _T_95532; // @[Mux.scala 31:69:@40388.4]
  wire [15:0] _T_95533; // @[Mux.scala 31:69:@40389.4]
  wire [15:0] _T_95534; // @[Mux.scala 31:69:@40390.4]
  wire [15:0] _T_95535; // @[Mux.scala 31:69:@40391.4]
  wire [15:0] _T_95536; // @[Mux.scala 31:69:@40392.4]
  wire [15:0] _T_95537; // @[Mux.scala 31:69:@40393.4]
  wire [15:0] _T_95538; // @[Mux.scala 31:69:@40394.4]
  wire [15:0] _T_95539; // @[Mux.scala 31:69:@40395.4]
  wire [15:0] _T_95540; // @[Mux.scala 31:69:@40396.4]
  wire [15:0] _T_95541; // @[Mux.scala 31:69:@40397.4]
  wire [15:0] _T_95542; // @[Mux.scala 31:69:@40398.4]
  wire  _T_95543; // @[OneHot.scala 66:30:@40399.4]
  wire  _T_95544; // @[OneHot.scala 66:30:@40400.4]
  wire  _T_95545; // @[OneHot.scala 66:30:@40401.4]
  wire  _T_95546; // @[OneHot.scala 66:30:@40402.4]
  wire  _T_95547; // @[OneHot.scala 66:30:@40403.4]
  wire  _T_95548; // @[OneHot.scala 66:30:@40404.4]
  wire  _T_95549; // @[OneHot.scala 66:30:@40405.4]
  wire  _T_95550; // @[OneHot.scala 66:30:@40406.4]
  wire  _T_95551; // @[OneHot.scala 66:30:@40407.4]
  wire  _T_95552; // @[OneHot.scala 66:30:@40408.4]
  wire  _T_95553; // @[OneHot.scala 66:30:@40409.4]
  wire  _T_95554; // @[OneHot.scala 66:30:@40410.4]
  wire  _T_95555; // @[OneHot.scala 66:30:@40411.4]
  wire  _T_95556; // @[OneHot.scala 66:30:@40412.4]
  wire  _T_95557; // @[OneHot.scala 66:30:@40413.4]
  wire  _T_95558; // @[OneHot.scala 66:30:@40414.4]
  wire [7:0] _T_95623; // @[Mux.scala 19:72:@40438.4]
  wire [15:0] _T_95631; // @[Mux.scala 19:72:@40446.4]
  wire [15:0] _T_95633; // @[Mux.scala 19:72:@40447.4]
  wire [7:0] _T_95640; // @[Mux.scala 19:72:@40454.4]
  wire [15:0] _T_95648; // @[Mux.scala 19:72:@40462.4]
  wire [15:0] _T_95650; // @[Mux.scala 19:72:@40463.4]
  wire [7:0] _T_95657; // @[Mux.scala 19:72:@40470.4]
  wire [15:0] _T_95665; // @[Mux.scala 19:72:@40478.4]
  wire [15:0] _T_95667; // @[Mux.scala 19:72:@40479.4]
  wire [7:0] _T_95674; // @[Mux.scala 19:72:@40486.4]
  wire [15:0] _T_95682; // @[Mux.scala 19:72:@40494.4]
  wire [15:0] _T_95684; // @[Mux.scala 19:72:@40495.4]
  wire [7:0] _T_95691; // @[Mux.scala 19:72:@40502.4]
  wire [15:0] _T_95699; // @[Mux.scala 19:72:@40510.4]
  wire [15:0] _T_95701; // @[Mux.scala 19:72:@40511.4]
  wire [7:0] _T_95708; // @[Mux.scala 19:72:@40518.4]
  wire [15:0] _T_95716; // @[Mux.scala 19:72:@40526.4]
  wire [15:0] _T_95718; // @[Mux.scala 19:72:@40527.4]
  wire [7:0] _T_95725; // @[Mux.scala 19:72:@40534.4]
  wire [15:0] _T_95733; // @[Mux.scala 19:72:@40542.4]
  wire [15:0] _T_95735; // @[Mux.scala 19:72:@40543.4]
  wire [7:0] _T_95742; // @[Mux.scala 19:72:@40550.4]
  wire [15:0] _T_95750; // @[Mux.scala 19:72:@40558.4]
  wire [15:0] _T_95752; // @[Mux.scala 19:72:@40559.4]
  wire [7:0] _T_95759; // @[Mux.scala 19:72:@40566.4]
  wire [15:0] _T_95767; // @[Mux.scala 19:72:@40574.4]
  wire [15:0] _T_95769; // @[Mux.scala 19:72:@40575.4]
  wire [7:0] _T_95776; // @[Mux.scala 19:72:@40582.4]
  wire [15:0] _T_95784; // @[Mux.scala 19:72:@40590.4]
  wire [15:0] _T_95786; // @[Mux.scala 19:72:@40591.4]
  wire [7:0] _T_95793; // @[Mux.scala 19:72:@40598.4]
  wire [15:0] _T_95801; // @[Mux.scala 19:72:@40606.4]
  wire [15:0] _T_95803; // @[Mux.scala 19:72:@40607.4]
  wire [7:0] _T_95810; // @[Mux.scala 19:72:@40614.4]
  wire [15:0] _T_95818; // @[Mux.scala 19:72:@40622.4]
  wire [15:0] _T_95820; // @[Mux.scala 19:72:@40623.4]
  wire [7:0] _T_95827; // @[Mux.scala 19:72:@40630.4]
  wire [15:0] _T_95835; // @[Mux.scala 19:72:@40638.4]
  wire [15:0] _T_95837; // @[Mux.scala 19:72:@40639.4]
  wire [7:0] _T_95844; // @[Mux.scala 19:72:@40646.4]
  wire [15:0] _T_95852; // @[Mux.scala 19:72:@40654.4]
  wire [15:0] _T_95854; // @[Mux.scala 19:72:@40655.4]
  wire [7:0] _T_95861; // @[Mux.scala 19:72:@40662.4]
  wire [15:0] _T_95869; // @[Mux.scala 19:72:@40670.4]
  wire [15:0] _T_95871; // @[Mux.scala 19:72:@40671.4]
  wire [7:0] _T_95878; // @[Mux.scala 19:72:@40678.4]
  wire [15:0] _T_95886; // @[Mux.scala 19:72:@40686.4]
  wire [15:0] _T_95888; // @[Mux.scala 19:72:@40687.4]
  wire [15:0] _T_95889; // @[Mux.scala 19:72:@40688.4]
  wire [15:0] _T_95890; // @[Mux.scala 19:72:@40689.4]
  wire [15:0] _T_95891; // @[Mux.scala 19:72:@40690.4]
  wire [15:0] _T_95892; // @[Mux.scala 19:72:@40691.4]
  wire [15:0] _T_95893; // @[Mux.scala 19:72:@40692.4]
  wire [15:0] _T_95894; // @[Mux.scala 19:72:@40693.4]
  wire [15:0] _T_95895; // @[Mux.scala 19:72:@40694.4]
  wire [15:0] _T_95896; // @[Mux.scala 19:72:@40695.4]
  wire [15:0] _T_95897; // @[Mux.scala 19:72:@40696.4]
  wire [15:0] _T_95898; // @[Mux.scala 19:72:@40697.4]
  wire [15:0] _T_95899; // @[Mux.scala 19:72:@40698.4]
  wire [15:0] _T_95900; // @[Mux.scala 19:72:@40699.4]
  wire [15:0] _T_95901; // @[Mux.scala 19:72:@40700.4]
  wire [15:0] _T_95902; // @[Mux.scala 19:72:@40701.4]
  wire [15:0] _T_95903; // @[Mux.scala 19:72:@40702.4]
  wire  inputPriorityPorts_0_0; // @[Mux.scala 19:72:@40706.4]
  wire  inputPriorityPorts_0_1; // @[Mux.scala 19:72:@40708.4]
  wire  inputPriorityPorts_0_2; // @[Mux.scala 19:72:@40710.4]
  wire  inputPriorityPorts_0_3; // @[Mux.scala 19:72:@40712.4]
  wire  inputPriorityPorts_0_4; // @[Mux.scala 19:72:@40714.4]
  wire  inputPriorityPorts_0_5; // @[Mux.scala 19:72:@40716.4]
  wire  inputPriorityPorts_0_6; // @[Mux.scala 19:72:@40718.4]
  wire  inputPriorityPorts_0_7; // @[Mux.scala 19:72:@40720.4]
  wire  inputPriorityPorts_0_8; // @[Mux.scala 19:72:@40722.4]
  wire  inputPriorityPorts_0_9; // @[Mux.scala 19:72:@40724.4]
  wire  inputPriorityPorts_0_10; // @[Mux.scala 19:72:@40726.4]
  wire  inputPriorityPorts_0_11; // @[Mux.scala 19:72:@40728.4]
  wire  inputPriorityPorts_0_12; // @[Mux.scala 19:72:@40730.4]
  wire  inputPriorityPorts_0_13; // @[Mux.scala 19:72:@40732.4]
  wire  inputPriorityPorts_0_14; // @[Mux.scala 19:72:@40734.4]
  wire  inputPriorityPorts_0_15; // @[Mux.scala 19:72:@40736.4]
  wire [15:0] _T_96105; // @[Mux.scala 31:69:@40790.4]
  wire [15:0] _T_96106; // @[Mux.scala 31:69:@40791.4]
  wire [15:0] _T_96107; // @[Mux.scala 31:69:@40792.4]
  wire [15:0] _T_96108; // @[Mux.scala 31:69:@40793.4]
  wire [15:0] _T_96109; // @[Mux.scala 31:69:@40794.4]
  wire [15:0] _T_96110; // @[Mux.scala 31:69:@40795.4]
  wire [15:0] _T_96111; // @[Mux.scala 31:69:@40796.4]
  wire [15:0] _T_96112; // @[Mux.scala 31:69:@40797.4]
  wire [15:0] _T_96113; // @[Mux.scala 31:69:@40798.4]
  wire [15:0] _T_96114; // @[Mux.scala 31:69:@40799.4]
  wire [15:0] _T_96115; // @[Mux.scala 31:69:@40800.4]
  wire [15:0] _T_96116; // @[Mux.scala 31:69:@40801.4]
  wire [15:0] _T_96117; // @[Mux.scala 31:69:@40802.4]
  wire [15:0] _T_96118; // @[Mux.scala 31:69:@40803.4]
  wire [15:0] _T_96119; // @[Mux.scala 31:69:@40804.4]
  wire [15:0] _T_96120; // @[Mux.scala 31:69:@40805.4]
  wire  _T_96121; // @[OneHot.scala 66:30:@40806.4]
  wire  _T_96122; // @[OneHot.scala 66:30:@40807.4]
  wire  _T_96123; // @[OneHot.scala 66:30:@40808.4]
  wire  _T_96124; // @[OneHot.scala 66:30:@40809.4]
  wire  _T_96125; // @[OneHot.scala 66:30:@40810.4]
  wire  _T_96126; // @[OneHot.scala 66:30:@40811.4]
  wire  _T_96127; // @[OneHot.scala 66:30:@40812.4]
  wire  _T_96128; // @[OneHot.scala 66:30:@40813.4]
  wire  _T_96129; // @[OneHot.scala 66:30:@40814.4]
  wire  _T_96130; // @[OneHot.scala 66:30:@40815.4]
  wire  _T_96131; // @[OneHot.scala 66:30:@40816.4]
  wire  _T_96132; // @[OneHot.scala 66:30:@40817.4]
  wire  _T_96133; // @[OneHot.scala 66:30:@40818.4]
  wire  _T_96134; // @[OneHot.scala 66:30:@40819.4]
  wire  _T_96135; // @[OneHot.scala 66:30:@40820.4]
  wire  _T_96136; // @[OneHot.scala 66:30:@40821.4]
  wire [15:0] _T_96177; // @[Mux.scala 31:69:@40839.4]
  wire [15:0] _T_96178; // @[Mux.scala 31:69:@40840.4]
  wire [15:0] _T_96179; // @[Mux.scala 31:69:@40841.4]
  wire [15:0] _T_96180; // @[Mux.scala 31:69:@40842.4]
  wire [15:0] _T_96181; // @[Mux.scala 31:69:@40843.4]
  wire [15:0] _T_96182; // @[Mux.scala 31:69:@40844.4]
  wire [15:0] _T_96183; // @[Mux.scala 31:69:@40845.4]
  wire [15:0] _T_96184; // @[Mux.scala 31:69:@40846.4]
  wire [15:0] _T_96185; // @[Mux.scala 31:69:@40847.4]
  wire [15:0] _T_96186; // @[Mux.scala 31:69:@40848.4]
  wire [15:0] _T_96187; // @[Mux.scala 31:69:@40849.4]
  wire [15:0] _T_96188; // @[Mux.scala 31:69:@40850.4]
  wire [15:0] _T_96189; // @[Mux.scala 31:69:@40851.4]
  wire [15:0] _T_96190; // @[Mux.scala 31:69:@40852.4]
  wire [15:0] _T_96191; // @[Mux.scala 31:69:@40853.4]
  wire [15:0] _T_96192; // @[Mux.scala 31:69:@40854.4]
  wire  _T_96193; // @[OneHot.scala 66:30:@40855.4]
  wire  _T_96194; // @[OneHot.scala 66:30:@40856.4]
  wire  _T_96195; // @[OneHot.scala 66:30:@40857.4]
  wire  _T_96196; // @[OneHot.scala 66:30:@40858.4]
  wire  _T_96197; // @[OneHot.scala 66:30:@40859.4]
  wire  _T_96198; // @[OneHot.scala 66:30:@40860.4]
  wire  _T_96199; // @[OneHot.scala 66:30:@40861.4]
  wire  _T_96200; // @[OneHot.scala 66:30:@40862.4]
  wire  _T_96201; // @[OneHot.scala 66:30:@40863.4]
  wire  _T_96202; // @[OneHot.scala 66:30:@40864.4]
  wire  _T_96203; // @[OneHot.scala 66:30:@40865.4]
  wire  _T_96204; // @[OneHot.scala 66:30:@40866.4]
  wire  _T_96205; // @[OneHot.scala 66:30:@40867.4]
  wire  _T_96206; // @[OneHot.scala 66:30:@40868.4]
  wire  _T_96207; // @[OneHot.scala 66:30:@40869.4]
  wire  _T_96208; // @[OneHot.scala 66:30:@40870.4]
  wire [15:0] _T_96249; // @[Mux.scala 31:69:@40888.4]
  wire [15:0] _T_96250; // @[Mux.scala 31:69:@40889.4]
  wire [15:0] _T_96251; // @[Mux.scala 31:69:@40890.4]
  wire [15:0] _T_96252; // @[Mux.scala 31:69:@40891.4]
  wire [15:0] _T_96253; // @[Mux.scala 31:69:@40892.4]
  wire [15:0] _T_96254; // @[Mux.scala 31:69:@40893.4]
  wire [15:0] _T_96255; // @[Mux.scala 31:69:@40894.4]
  wire [15:0] _T_96256; // @[Mux.scala 31:69:@40895.4]
  wire [15:0] _T_96257; // @[Mux.scala 31:69:@40896.4]
  wire [15:0] _T_96258; // @[Mux.scala 31:69:@40897.4]
  wire [15:0] _T_96259; // @[Mux.scala 31:69:@40898.4]
  wire [15:0] _T_96260; // @[Mux.scala 31:69:@40899.4]
  wire [15:0] _T_96261; // @[Mux.scala 31:69:@40900.4]
  wire [15:0] _T_96262; // @[Mux.scala 31:69:@40901.4]
  wire [15:0] _T_96263; // @[Mux.scala 31:69:@40902.4]
  wire [15:0] _T_96264; // @[Mux.scala 31:69:@40903.4]
  wire  _T_96265; // @[OneHot.scala 66:30:@40904.4]
  wire  _T_96266; // @[OneHot.scala 66:30:@40905.4]
  wire  _T_96267; // @[OneHot.scala 66:30:@40906.4]
  wire  _T_96268; // @[OneHot.scala 66:30:@40907.4]
  wire  _T_96269; // @[OneHot.scala 66:30:@40908.4]
  wire  _T_96270; // @[OneHot.scala 66:30:@40909.4]
  wire  _T_96271; // @[OneHot.scala 66:30:@40910.4]
  wire  _T_96272; // @[OneHot.scala 66:30:@40911.4]
  wire  _T_96273; // @[OneHot.scala 66:30:@40912.4]
  wire  _T_96274; // @[OneHot.scala 66:30:@40913.4]
  wire  _T_96275; // @[OneHot.scala 66:30:@40914.4]
  wire  _T_96276; // @[OneHot.scala 66:30:@40915.4]
  wire  _T_96277; // @[OneHot.scala 66:30:@40916.4]
  wire  _T_96278; // @[OneHot.scala 66:30:@40917.4]
  wire  _T_96279; // @[OneHot.scala 66:30:@40918.4]
  wire  _T_96280; // @[OneHot.scala 66:30:@40919.4]
  wire [15:0] _T_96321; // @[Mux.scala 31:69:@40937.4]
  wire [15:0] _T_96322; // @[Mux.scala 31:69:@40938.4]
  wire [15:0] _T_96323; // @[Mux.scala 31:69:@40939.4]
  wire [15:0] _T_96324; // @[Mux.scala 31:69:@40940.4]
  wire [15:0] _T_96325; // @[Mux.scala 31:69:@40941.4]
  wire [15:0] _T_96326; // @[Mux.scala 31:69:@40942.4]
  wire [15:0] _T_96327; // @[Mux.scala 31:69:@40943.4]
  wire [15:0] _T_96328; // @[Mux.scala 31:69:@40944.4]
  wire [15:0] _T_96329; // @[Mux.scala 31:69:@40945.4]
  wire [15:0] _T_96330; // @[Mux.scala 31:69:@40946.4]
  wire [15:0] _T_96331; // @[Mux.scala 31:69:@40947.4]
  wire [15:0] _T_96332; // @[Mux.scala 31:69:@40948.4]
  wire [15:0] _T_96333; // @[Mux.scala 31:69:@40949.4]
  wire [15:0] _T_96334; // @[Mux.scala 31:69:@40950.4]
  wire [15:0] _T_96335; // @[Mux.scala 31:69:@40951.4]
  wire [15:0] _T_96336; // @[Mux.scala 31:69:@40952.4]
  wire  _T_96337; // @[OneHot.scala 66:30:@40953.4]
  wire  _T_96338; // @[OneHot.scala 66:30:@40954.4]
  wire  _T_96339; // @[OneHot.scala 66:30:@40955.4]
  wire  _T_96340; // @[OneHot.scala 66:30:@40956.4]
  wire  _T_96341; // @[OneHot.scala 66:30:@40957.4]
  wire  _T_96342; // @[OneHot.scala 66:30:@40958.4]
  wire  _T_96343; // @[OneHot.scala 66:30:@40959.4]
  wire  _T_96344; // @[OneHot.scala 66:30:@40960.4]
  wire  _T_96345; // @[OneHot.scala 66:30:@40961.4]
  wire  _T_96346; // @[OneHot.scala 66:30:@40962.4]
  wire  _T_96347; // @[OneHot.scala 66:30:@40963.4]
  wire  _T_96348; // @[OneHot.scala 66:30:@40964.4]
  wire  _T_96349; // @[OneHot.scala 66:30:@40965.4]
  wire  _T_96350; // @[OneHot.scala 66:30:@40966.4]
  wire  _T_96351; // @[OneHot.scala 66:30:@40967.4]
  wire  _T_96352; // @[OneHot.scala 66:30:@40968.4]
  wire [15:0] _T_96393; // @[Mux.scala 31:69:@40986.4]
  wire [15:0] _T_96394; // @[Mux.scala 31:69:@40987.4]
  wire [15:0] _T_96395; // @[Mux.scala 31:69:@40988.4]
  wire [15:0] _T_96396; // @[Mux.scala 31:69:@40989.4]
  wire [15:0] _T_96397; // @[Mux.scala 31:69:@40990.4]
  wire [15:0] _T_96398; // @[Mux.scala 31:69:@40991.4]
  wire [15:0] _T_96399; // @[Mux.scala 31:69:@40992.4]
  wire [15:0] _T_96400; // @[Mux.scala 31:69:@40993.4]
  wire [15:0] _T_96401; // @[Mux.scala 31:69:@40994.4]
  wire [15:0] _T_96402; // @[Mux.scala 31:69:@40995.4]
  wire [15:0] _T_96403; // @[Mux.scala 31:69:@40996.4]
  wire [15:0] _T_96404; // @[Mux.scala 31:69:@40997.4]
  wire [15:0] _T_96405; // @[Mux.scala 31:69:@40998.4]
  wire [15:0] _T_96406; // @[Mux.scala 31:69:@40999.4]
  wire [15:0] _T_96407; // @[Mux.scala 31:69:@41000.4]
  wire [15:0] _T_96408; // @[Mux.scala 31:69:@41001.4]
  wire  _T_96409; // @[OneHot.scala 66:30:@41002.4]
  wire  _T_96410; // @[OneHot.scala 66:30:@41003.4]
  wire  _T_96411; // @[OneHot.scala 66:30:@41004.4]
  wire  _T_96412; // @[OneHot.scala 66:30:@41005.4]
  wire  _T_96413; // @[OneHot.scala 66:30:@41006.4]
  wire  _T_96414; // @[OneHot.scala 66:30:@41007.4]
  wire  _T_96415; // @[OneHot.scala 66:30:@41008.4]
  wire  _T_96416; // @[OneHot.scala 66:30:@41009.4]
  wire  _T_96417; // @[OneHot.scala 66:30:@41010.4]
  wire  _T_96418; // @[OneHot.scala 66:30:@41011.4]
  wire  _T_96419; // @[OneHot.scala 66:30:@41012.4]
  wire  _T_96420; // @[OneHot.scala 66:30:@41013.4]
  wire  _T_96421; // @[OneHot.scala 66:30:@41014.4]
  wire  _T_96422; // @[OneHot.scala 66:30:@41015.4]
  wire  _T_96423; // @[OneHot.scala 66:30:@41016.4]
  wire  _T_96424; // @[OneHot.scala 66:30:@41017.4]
  wire [15:0] _T_96465; // @[Mux.scala 31:69:@41035.4]
  wire [15:0] _T_96466; // @[Mux.scala 31:69:@41036.4]
  wire [15:0] _T_96467; // @[Mux.scala 31:69:@41037.4]
  wire [15:0] _T_96468; // @[Mux.scala 31:69:@41038.4]
  wire [15:0] _T_96469; // @[Mux.scala 31:69:@41039.4]
  wire [15:0] _T_96470; // @[Mux.scala 31:69:@41040.4]
  wire [15:0] _T_96471; // @[Mux.scala 31:69:@41041.4]
  wire [15:0] _T_96472; // @[Mux.scala 31:69:@41042.4]
  wire [15:0] _T_96473; // @[Mux.scala 31:69:@41043.4]
  wire [15:0] _T_96474; // @[Mux.scala 31:69:@41044.4]
  wire [15:0] _T_96475; // @[Mux.scala 31:69:@41045.4]
  wire [15:0] _T_96476; // @[Mux.scala 31:69:@41046.4]
  wire [15:0] _T_96477; // @[Mux.scala 31:69:@41047.4]
  wire [15:0] _T_96478; // @[Mux.scala 31:69:@41048.4]
  wire [15:0] _T_96479; // @[Mux.scala 31:69:@41049.4]
  wire [15:0] _T_96480; // @[Mux.scala 31:69:@41050.4]
  wire  _T_96481; // @[OneHot.scala 66:30:@41051.4]
  wire  _T_96482; // @[OneHot.scala 66:30:@41052.4]
  wire  _T_96483; // @[OneHot.scala 66:30:@41053.4]
  wire  _T_96484; // @[OneHot.scala 66:30:@41054.4]
  wire  _T_96485; // @[OneHot.scala 66:30:@41055.4]
  wire  _T_96486; // @[OneHot.scala 66:30:@41056.4]
  wire  _T_96487; // @[OneHot.scala 66:30:@41057.4]
  wire  _T_96488; // @[OneHot.scala 66:30:@41058.4]
  wire  _T_96489; // @[OneHot.scala 66:30:@41059.4]
  wire  _T_96490; // @[OneHot.scala 66:30:@41060.4]
  wire  _T_96491; // @[OneHot.scala 66:30:@41061.4]
  wire  _T_96492; // @[OneHot.scala 66:30:@41062.4]
  wire  _T_96493; // @[OneHot.scala 66:30:@41063.4]
  wire  _T_96494; // @[OneHot.scala 66:30:@41064.4]
  wire  _T_96495; // @[OneHot.scala 66:30:@41065.4]
  wire  _T_96496; // @[OneHot.scala 66:30:@41066.4]
  wire [15:0] _T_96537; // @[Mux.scala 31:69:@41084.4]
  wire [15:0] _T_96538; // @[Mux.scala 31:69:@41085.4]
  wire [15:0] _T_96539; // @[Mux.scala 31:69:@41086.4]
  wire [15:0] _T_96540; // @[Mux.scala 31:69:@41087.4]
  wire [15:0] _T_96541; // @[Mux.scala 31:69:@41088.4]
  wire [15:0] _T_96542; // @[Mux.scala 31:69:@41089.4]
  wire [15:0] _T_96543; // @[Mux.scala 31:69:@41090.4]
  wire [15:0] _T_96544; // @[Mux.scala 31:69:@41091.4]
  wire [15:0] _T_96545; // @[Mux.scala 31:69:@41092.4]
  wire [15:0] _T_96546; // @[Mux.scala 31:69:@41093.4]
  wire [15:0] _T_96547; // @[Mux.scala 31:69:@41094.4]
  wire [15:0] _T_96548; // @[Mux.scala 31:69:@41095.4]
  wire [15:0] _T_96549; // @[Mux.scala 31:69:@41096.4]
  wire [15:0] _T_96550; // @[Mux.scala 31:69:@41097.4]
  wire [15:0] _T_96551; // @[Mux.scala 31:69:@41098.4]
  wire [15:0] _T_96552; // @[Mux.scala 31:69:@41099.4]
  wire  _T_96553; // @[OneHot.scala 66:30:@41100.4]
  wire  _T_96554; // @[OneHot.scala 66:30:@41101.4]
  wire  _T_96555; // @[OneHot.scala 66:30:@41102.4]
  wire  _T_96556; // @[OneHot.scala 66:30:@41103.4]
  wire  _T_96557; // @[OneHot.scala 66:30:@41104.4]
  wire  _T_96558; // @[OneHot.scala 66:30:@41105.4]
  wire  _T_96559; // @[OneHot.scala 66:30:@41106.4]
  wire  _T_96560; // @[OneHot.scala 66:30:@41107.4]
  wire  _T_96561; // @[OneHot.scala 66:30:@41108.4]
  wire  _T_96562; // @[OneHot.scala 66:30:@41109.4]
  wire  _T_96563; // @[OneHot.scala 66:30:@41110.4]
  wire  _T_96564; // @[OneHot.scala 66:30:@41111.4]
  wire  _T_96565; // @[OneHot.scala 66:30:@41112.4]
  wire  _T_96566; // @[OneHot.scala 66:30:@41113.4]
  wire  _T_96567; // @[OneHot.scala 66:30:@41114.4]
  wire  _T_96568; // @[OneHot.scala 66:30:@41115.4]
  wire [15:0] _T_96609; // @[Mux.scala 31:69:@41133.4]
  wire [15:0] _T_96610; // @[Mux.scala 31:69:@41134.4]
  wire [15:0] _T_96611; // @[Mux.scala 31:69:@41135.4]
  wire [15:0] _T_96612; // @[Mux.scala 31:69:@41136.4]
  wire [15:0] _T_96613; // @[Mux.scala 31:69:@41137.4]
  wire [15:0] _T_96614; // @[Mux.scala 31:69:@41138.4]
  wire [15:0] _T_96615; // @[Mux.scala 31:69:@41139.4]
  wire [15:0] _T_96616; // @[Mux.scala 31:69:@41140.4]
  wire [15:0] _T_96617; // @[Mux.scala 31:69:@41141.4]
  wire [15:0] _T_96618; // @[Mux.scala 31:69:@41142.4]
  wire [15:0] _T_96619; // @[Mux.scala 31:69:@41143.4]
  wire [15:0] _T_96620; // @[Mux.scala 31:69:@41144.4]
  wire [15:0] _T_96621; // @[Mux.scala 31:69:@41145.4]
  wire [15:0] _T_96622; // @[Mux.scala 31:69:@41146.4]
  wire [15:0] _T_96623; // @[Mux.scala 31:69:@41147.4]
  wire [15:0] _T_96624; // @[Mux.scala 31:69:@41148.4]
  wire  _T_96625; // @[OneHot.scala 66:30:@41149.4]
  wire  _T_96626; // @[OneHot.scala 66:30:@41150.4]
  wire  _T_96627; // @[OneHot.scala 66:30:@41151.4]
  wire  _T_96628; // @[OneHot.scala 66:30:@41152.4]
  wire  _T_96629; // @[OneHot.scala 66:30:@41153.4]
  wire  _T_96630; // @[OneHot.scala 66:30:@41154.4]
  wire  _T_96631; // @[OneHot.scala 66:30:@41155.4]
  wire  _T_96632; // @[OneHot.scala 66:30:@41156.4]
  wire  _T_96633; // @[OneHot.scala 66:30:@41157.4]
  wire  _T_96634; // @[OneHot.scala 66:30:@41158.4]
  wire  _T_96635; // @[OneHot.scala 66:30:@41159.4]
  wire  _T_96636; // @[OneHot.scala 66:30:@41160.4]
  wire  _T_96637; // @[OneHot.scala 66:30:@41161.4]
  wire  _T_96638; // @[OneHot.scala 66:30:@41162.4]
  wire  _T_96639; // @[OneHot.scala 66:30:@41163.4]
  wire  _T_96640; // @[OneHot.scala 66:30:@41164.4]
  wire [15:0] _T_96681; // @[Mux.scala 31:69:@41182.4]
  wire [15:0] _T_96682; // @[Mux.scala 31:69:@41183.4]
  wire [15:0] _T_96683; // @[Mux.scala 31:69:@41184.4]
  wire [15:0] _T_96684; // @[Mux.scala 31:69:@41185.4]
  wire [15:0] _T_96685; // @[Mux.scala 31:69:@41186.4]
  wire [15:0] _T_96686; // @[Mux.scala 31:69:@41187.4]
  wire [15:0] _T_96687; // @[Mux.scala 31:69:@41188.4]
  wire [15:0] _T_96688; // @[Mux.scala 31:69:@41189.4]
  wire [15:0] _T_96689; // @[Mux.scala 31:69:@41190.4]
  wire [15:0] _T_96690; // @[Mux.scala 31:69:@41191.4]
  wire [15:0] _T_96691; // @[Mux.scala 31:69:@41192.4]
  wire [15:0] _T_96692; // @[Mux.scala 31:69:@41193.4]
  wire [15:0] _T_96693; // @[Mux.scala 31:69:@41194.4]
  wire [15:0] _T_96694; // @[Mux.scala 31:69:@41195.4]
  wire [15:0] _T_96695; // @[Mux.scala 31:69:@41196.4]
  wire [15:0] _T_96696; // @[Mux.scala 31:69:@41197.4]
  wire  _T_96697; // @[OneHot.scala 66:30:@41198.4]
  wire  _T_96698; // @[OneHot.scala 66:30:@41199.4]
  wire  _T_96699; // @[OneHot.scala 66:30:@41200.4]
  wire  _T_96700; // @[OneHot.scala 66:30:@41201.4]
  wire  _T_96701; // @[OneHot.scala 66:30:@41202.4]
  wire  _T_96702; // @[OneHot.scala 66:30:@41203.4]
  wire  _T_96703; // @[OneHot.scala 66:30:@41204.4]
  wire  _T_96704; // @[OneHot.scala 66:30:@41205.4]
  wire  _T_96705; // @[OneHot.scala 66:30:@41206.4]
  wire  _T_96706; // @[OneHot.scala 66:30:@41207.4]
  wire  _T_96707; // @[OneHot.scala 66:30:@41208.4]
  wire  _T_96708; // @[OneHot.scala 66:30:@41209.4]
  wire  _T_96709; // @[OneHot.scala 66:30:@41210.4]
  wire  _T_96710; // @[OneHot.scala 66:30:@41211.4]
  wire  _T_96711; // @[OneHot.scala 66:30:@41212.4]
  wire  _T_96712; // @[OneHot.scala 66:30:@41213.4]
  wire [15:0] _T_96753; // @[Mux.scala 31:69:@41231.4]
  wire [15:0] _T_96754; // @[Mux.scala 31:69:@41232.4]
  wire [15:0] _T_96755; // @[Mux.scala 31:69:@41233.4]
  wire [15:0] _T_96756; // @[Mux.scala 31:69:@41234.4]
  wire [15:0] _T_96757; // @[Mux.scala 31:69:@41235.4]
  wire [15:0] _T_96758; // @[Mux.scala 31:69:@41236.4]
  wire [15:0] _T_96759; // @[Mux.scala 31:69:@41237.4]
  wire [15:0] _T_96760; // @[Mux.scala 31:69:@41238.4]
  wire [15:0] _T_96761; // @[Mux.scala 31:69:@41239.4]
  wire [15:0] _T_96762; // @[Mux.scala 31:69:@41240.4]
  wire [15:0] _T_96763; // @[Mux.scala 31:69:@41241.4]
  wire [15:0] _T_96764; // @[Mux.scala 31:69:@41242.4]
  wire [15:0] _T_96765; // @[Mux.scala 31:69:@41243.4]
  wire [15:0] _T_96766; // @[Mux.scala 31:69:@41244.4]
  wire [15:0] _T_96767; // @[Mux.scala 31:69:@41245.4]
  wire [15:0] _T_96768; // @[Mux.scala 31:69:@41246.4]
  wire  _T_96769; // @[OneHot.scala 66:30:@41247.4]
  wire  _T_96770; // @[OneHot.scala 66:30:@41248.4]
  wire  _T_96771; // @[OneHot.scala 66:30:@41249.4]
  wire  _T_96772; // @[OneHot.scala 66:30:@41250.4]
  wire  _T_96773; // @[OneHot.scala 66:30:@41251.4]
  wire  _T_96774; // @[OneHot.scala 66:30:@41252.4]
  wire  _T_96775; // @[OneHot.scala 66:30:@41253.4]
  wire  _T_96776; // @[OneHot.scala 66:30:@41254.4]
  wire  _T_96777; // @[OneHot.scala 66:30:@41255.4]
  wire  _T_96778; // @[OneHot.scala 66:30:@41256.4]
  wire  _T_96779; // @[OneHot.scala 66:30:@41257.4]
  wire  _T_96780; // @[OneHot.scala 66:30:@41258.4]
  wire  _T_96781; // @[OneHot.scala 66:30:@41259.4]
  wire  _T_96782; // @[OneHot.scala 66:30:@41260.4]
  wire  _T_96783; // @[OneHot.scala 66:30:@41261.4]
  wire  _T_96784; // @[OneHot.scala 66:30:@41262.4]
  wire [15:0] _T_96825; // @[Mux.scala 31:69:@41280.4]
  wire [15:0] _T_96826; // @[Mux.scala 31:69:@41281.4]
  wire [15:0] _T_96827; // @[Mux.scala 31:69:@41282.4]
  wire [15:0] _T_96828; // @[Mux.scala 31:69:@41283.4]
  wire [15:0] _T_96829; // @[Mux.scala 31:69:@41284.4]
  wire [15:0] _T_96830; // @[Mux.scala 31:69:@41285.4]
  wire [15:0] _T_96831; // @[Mux.scala 31:69:@41286.4]
  wire [15:0] _T_96832; // @[Mux.scala 31:69:@41287.4]
  wire [15:0] _T_96833; // @[Mux.scala 31:69:@41288.4]
  wire [15:0] _T_96834; // @[Mux.scala 31:69:@41289.4]
  wire [15:0] _T_96835; // @[Mux.scala 31:69:@41290.4]
  wire [15:0] _T_96836; // @[Mux.scala 31:69:@41291.4]
  wire [15:0] _T_96837; // @[Mux.scala 31:69:@41292.4]
  wire [15:0] _T_96838; // @[Mux.scala 31:69:@41293.4]
  wire [15:0] _T_96839; // @[Mux.scala 31:69:@41294.4]
  wire [15:0] _T_96840; // @[Mux.scala 31:69:@41295.4]
  wire  _T_96841; // @[OneHot.scala 66:30:@41296.4]
  wire  _T_96842; // @[OneHot.scala 66:30:@41297.4]
  wire  _T_96843; // @[OneHot.scala 66:30:@41298.4]
  wire  _T_96844; // @[OneHot.scala 66:30:@41299.4]
  wire  _T_96845; // @[OneHot.scala 66:30:@41300.4]
  wire  _T_96846; // @[OneHot.scala 66:30:@41301.4]
  wire  _T_96847; // @[OneHot.scala 66:30:@41302.4]
  wire  _T_96848; // @[OneHot.scala 66:30:@41303.4]
  wire  _T_96849; // @[OneHot.scala 66:30:@41304.4]
  wire  _T_96850; // @[OneHot.scala 66:30:@41305.4]
  wire  _T_96851; // @[OneHot.scala 66:30:@41306.4]
  wire  _T_96852; // @[OneHot.scala 66:30:@41307.4]
  wire  _T_96853; // @[OneHot.scala 66:30:@41308.4]
  wire  _T_96854; // @[OneHot.scala 66:30:@41309.4]
  wire  _T_96855; // @[OneHot.scala 66:30:@41310.4]
  wire  _T_96856; // @[OneHot.scala 66:30:@41311.4]
  wire [15:0] _T_96897; // @[Mux.scala 31:69:@41329.4]
  wire [15:0] _T_96898; // @[Mux.scala 31:69:@41330.4]
  wire [15:0] _T_96899; // @[Mux.scala 31:69:@41331.4]
  wire [15:0] _T_96900; // @[Mux.scala 31:69:@41332.4]
  wire [15:0] _T_96901; // @[Mux.scala 31:69:@41333.4]
  wire [15:0] _T_96902; // @[Mux.scala 31:69:@41334.4]
  wire [15:0] _T_96903; // @[Mux.scala 31:69:@41335.4]
  wire [15:0] _T_96904; // @[Mux.scala 31:69:@41336.4]
  wire [15:0] _T_96905; // @[Mux.scala 31:69:@41337.4]
  wire [15:0] _T_96906; // @[Mux.scala 31:69:@41338.4]
  wire [15:0] _T_96907; // @[Mux.scala 31:69:@41339.4]
  wire [15:0] _T_96908; // @[Mux.scala 31:69:@41340.4]
  wire [15:0] _T_96909; // @[Mux.scala 31:69:@41341.4]
  wire [15:0] _T_96910; // @[Mux.scala 31:69:@41342.4]
  wire [15:0] _T_96911; // @[Mux.scala 31:69:@41343.4]
  wire [15:0] _T_96912; // @[Mux.scala 31:69:@41344.4]
  wire  _T_96913; // @[OneHot.scala 66:30:@41345.4]
  wire  _T_96914; // @[OneHot.scala 66:30:@41346.4]
  wire  _T_96915; // @[OneHot.scala 66:30:@41347.4]
  wire  _T_96916; // @[OneHot.scala 66:30:@41348.4]
  wire  _T_96917; // @[OneHot.scala 66:30:@41349.4]
  wire  _T_96918; // @[OneHot.scala 66:30:@41350.4]
  wire  _T_96919; // @[OneHot.scala 66:30:@41351.4]
  wire  _T_96920; // @[OneHot.scala 66:30:@41352.4]
  wire  _T_96921; // @[OneHot.scala 66:30:@41353.4]
  wire  _T_96922; // @[OneHot.scala 66:30:@41354.4]
  wire  _T_96923; // @[OneHot.scala 66:30:@41355.4]
  wire  _T_96924; // @[OneHot.scala 66:30:@41356.4]
  wire  _T_96925; // @[OneHot.scala 66:30:@41357.4]
  wire  _T_96926; // @[OneHot.scala 66:30:@41358.4]
  wire  _T_96927; // @[OneHot.scala 66:30:@41359.4]
  wire  _T_96928; // @[OneHot.scala 66:30:@41360.4]
  wire [15:0] _T_96969; // @[Mux.scala 31:69:@41378.4]
  wire [15:0] _T_96970; // @[Mux.scala 31:69:@41379.4]
  wire [15:0] _T_96971; // @[Mux.scala 31:69:@41380.4]
  wire [15:0] _T_96972; // @[Mux.scala 31:69:@41381.4]
  wire [15:0] _T_96973; // @[Mux.scala 31:69:@41382.4]
  wire [15:0] _T_96974; // @[Mux.scala 31:69:@41383.4]
  wire [15:0] _T_96975; // @[Mux.scala 31:69:@41384.4]
  wire [15:0] _T_96976; // @[Mux.scala 31:69:@41385.4]
  wire [15:0] _T_96977; // @[Mux.scala 31:69:@41386.4]
  wire [15:0] _T_96978; // @[Mux.scala 31:69:@41387.4]
  wire [15:0] _T_96979; // @[Mux.scala 31:69:@41388.4]
  wire [15:0] _T_96980; // @[Mux.scala 31:69:@41389.4]
  wire [15:0] _T_96981; // @[Mux.scala 31:69:@41390.4]
  wire [15:0] _T_96982; // @[Mux.scala 31:69:@41391.4]
  wire [15:0] _T_96983; // @[Mux.scala 31:69:@41392.4]
  wire [15:0] _T_96984; // @[Mux.scala 31:69:@41393.4]
  wire  _T_96985; // @[OneHot.scala 66:30:@41394.4]
  wire  _T_96986; // @[OneHot.scala 66:30:@41395.4]
  wire  _T_96987; // @[OneHot.scala 66:30:@41396.4]
  wire  _T_96988; // @[OneHot.scala 66:30:@41397.4]
  wire  _T_96989; // @[OneHot.scala 66:30:@41398.4]
  wire  _T_96990; // @[OneHot.scala 66:30:@41399.4]
  wire  _T_96991; // @[OneHot.scala 66:30:@41400.4]
  wire  _T_96992; // @[OneHot.scala 66:30:@41401.4]
  wire  _T_96993; // @[OneHot.scala 66:30:@41402.4]
  wire  _T_96994; // @[OneHot.scala 66:30:@41403.4]
  wire  _T_96995; // @[OneHot.scala 66:30:@41404.4]
  wire  _T_96996; // @[OneHot.scala 66:30:@41405.4]
  wire  _T_96997; // @[OneHot.scala 66:30:@41406.4]
  wire  _T_96998; // @[OneHot.scala 66:30:@41407.4]
  wire  _T_96999; // @[OneHot.scala 66:30:@41408.4]
  wire  _T_97000; // @[OneHot.scala 66:30:@41409.4]
  wire [15:0] _T_97041; // @[Mux.scala 31:69:@41427.4]
  wire [15:0] _T_97042; // @[Mux.scala 31:69:@41428.4]
  wire [15:0] _T_97043; // @[Mux.scala 31:69:@41429.4]
  wire [15:0] _T_97044; // @[Mux.scala 31:69:@41430.4]
  wire [15:0] _T_97045; // @[Mux.scala 31:69:@41431.4]
  wire [15:0] _T_97046; // @[Mux.scala 31:69:@41432.4]
  wire [15:0] _T_97047; // @[Mux.scala 31:69:@41433.4]
  wire [15:0] _T_97048; // @[Mux.scala 31:69:@41434.4]
  wire [15:0] _T_97049; // @[Mux.scala 31:69:@41435.4]
  wire [15:0] _T_97050; // @[Mux.scala 31:69:@41436.4]
  wire [15:0] _T_97051; // @[Mux.scala 31:69:@41437.4]
  wire [15:0] _T_97052; // @[Mux.scala 31:69:@41438.4]
  wire [15:0] _T_97053; // @[Mux.scala 31:69:@41439.4]
  wire [15:0] _T_97054; // @[Mux.scala 31:69:@41440.4]
  wire [15:0] _T_97055; // @[Mux.scala 31:69:@41441.4]
  wire [15:0] _T_97056; // @[Mux.scala 31:69:@41442.4]
  wire  _T_97057; // @[OneHot.scala 66:30:@41443.4]
  wire  _T_97058; // @[OneHot.scala 66:30:@41444.4]
  wire  _T_97059; // @[OneHot.scala 66:30:@41445.4]
  wire  _T_97060; // @[OneHot.scala 66:30:@41446.4]
  wire  _T_97061; // @[OneHot.scala 66:30:@41447.4]
  wire  _T_97062; // @[OneHot.scala 66:30:@41448.4]
  wire  _T_97063; // @[OneHot.scala 66:30:@41449.4]
  wire  _T_97064; // @[OneHot.scala 66:30:@41450.4]
  wire  _T_97065; // @[OneHot.scala 66:30:@41451.4]
  wire  _T_97066; // @[OneHot.scala 66:30:@41452.4]
  wire  _T_97067; // @[OneHot.scala 66:30:@41453.4]
  wire  _T_97068; // @[OneHot.scala 66:30:@41454.4]
  wire  _T_97069; // @[OneHot.scala 66:30:@41455.4]
  wire  _T_97070; // @[OneHot.scala 66:30:@41456.4]
  wire  _T_97071; // @[OneHot.scala 66:30:@41457.4]
  wire  _T_97072; // @[OneHot.scala 66:30:@41458.4]
  wire [15:0] _T_97113; // @[Mux.scala 31:69:@41476.4]
  wire [15:0] _T_97114; // @[Mux.scala 31:69:@41477.4]
  wire [15:0] _T_97115; // @[Mux.scala 31:69:@41478.4]
  wire [15:0] _T_97116; // @[Mux.scala 31:69:@41479.4]
  wire [15:0] _T_97117; // @[Mux.scala 31:69:@41480.4]
  wire [15:0] _T_97118; // @[Mux.scala 31:69:@41481.4]
  wire [15:0] _T_97119; // @[Mux.scala 31:69:@41482.4]
  wire [15:0] _T_97120; // @[Mux.scala 31:69:@41483.4]
  wire [15:0] _T_97121; // @[Mux.scala 31:69:@41484.4]
  wire [15:0] _T_97122; // @[Mux.scala 31:69:@41485.4]
  wire [15:0] _T_97123; // @[Mux.scala 31:69:@41486.4]
  wire [15:0] _T_97124; // @[Mux.scala 31:69:@41487.4]
  wire [15:0] _T_97125; // @[Mux.scala 31:69:@41488.4]
  wire [15:0] _T_97126; // @[Mux.scala 31:69:@41489.4]
  wire [15:0] _T_97127; // @[Mux.scala 31:69:@41490.4]
  wire [15:0] _T_97128; // @[Mux.scala 31:69:@41491.4]
  wire  _T_97129; // @[OneHot.scala 66:30:@41492.4]
  wire  _T_97130; // @[OneHot.scala 66:30:@41493.4]
  wire  _T_97131; // @[OneHot.scala 66:30:@41494.4]
  wire  _T_97132; // @[OneHot.scala 66:30:@41495.4]
  wire  _T_97133; // @[OneHot.scala 66:30:@41496.4]
  wire  _T_97134; // @[OneHot.scala 66:30:@41497.4]
  wire  _T_97135; // @[OneHot.scala 66:30:@41498.4]
  wire  _T_97136; // @[OneHot.scala 66:30:@41499.4]
  wire  _T_97137; // @[OneHot.scala 66:30:@41500.4]
  wire  _T_97138; // @[OneHot.scala 66:30:@41501.4]
  wire  _T_97139; // @[OneHot.scala 66:30:@41502.4]
  wire  _T_97140; // @[OneHot.scala 66:30:@41503.4]
  wire  _T_97141; // @[OneHot.scala 66:30:@41504.4]
  wire  _T_97142; // @[OneHot.scala 66:30:@41505.4]
  wire  _T_97143; // @[OneHot.scala 66:30:@41506.4]
  wire  _T_97144; // @[OneHot.scala 66:30:@41507.4]
  wire [15:0] _T_97185; // @[Mux.scala 31:69:@41525.4]
  wire [15:0] _T_97186; // @[Mux.scala 31:69:@41526.4]
  wire [15:0] _T_97187; // @[Mux.scala 31:69:@41527.4]
  wire [15:0] _T_97188; // @[Mux.scala 31:69:@41528.4]
  wire [15:0] _T_97189; // @[Mux.scala 31:69:@41529.4]
  wire [15:0] _T_97190; // @[Mux.scala 31:69:@41530.4]
  wire [15:0] _T_97191; // @[Mux.scala 31:69:@41531.4]
  wire [15:0] _T_97192; // @[Mux.scala 31:69:@41532.4]
  wire [15:0] _T_97193; // @[Mux.scala 31:69:@41533.4]
  wire [15:0] _T_97194; // @[Mux.scala 31:69:@41534.4]
  wire [15:0] _T_97195; // @[Mux.scala 31:69:@41535.4]
  wire [15:0] _T_97196; // @[Mux.scala 31:69:@41536.4]
  wire [15:0] _T_97197; // @[Mux.scala 31:69:@41537.4]
  wire [15:0] _T_97198; // @[Mux.scala 31:69:@41538.4]
  wire [15:0] _T_97199; // @[Mux.scala 31:69:@41539.4]
  wire [15:0] _T_97200; // @[Mux.scala 31:69:@41540.4]
  wire  _T_97201; // @[OneHot.scala 66:30:@41541.4]
  wire  _T_97202; // @[OneHot.scala 66:30:@41542.4]
  wire  _T_97203; // @[OneHot.scala 66:30:@41543.4]
  wire  _T_97204; // @[OneHot.scala 66:30:@41544.4]
  wire  _T_97205; // @[OneHot.scala 66:30:@41545.4]
  wire  _T_97206; // @[OneHot.scala 66:30:@41546.4]
  wire  _T_97207; // @[OneHot.scala 66:30:@41547.4]
  wire  _T_97208; // @[OneHot.scala 66:30:@41548.4]
  wire  _T_97209; // @[OneHot.scala 66:30:@41549.4]
  wire  _T_97210; // @[OneHot.scala 66:30:@41550.4]
  wire  _T_97211; // @[OneHot.scala 66:30:@41551.4]
  wire  _T_97212; // @[OneHot.scala 66:30:@41552.4]
  wire  _T_97213; // @[OneHot.scala 66:30:@41553.4]
  wire  _T_97214; // @[OneHot.scala 66:30:@41554.4]
  wire  _T_97215; // @[OneHot.scala 66:30:@41555.4]
  wire  _T_97216; // @[OneHot.scala 66:30:@41556.4]
  wire [7:0] _T_97281; // @[Mux.scala 19:72:@41580.4]
  wire [15:0] _T_97289; // @[Mux.scala 19:72:@41588.4]
  wire [15:0] _T_97291; // @[Mux.scala 19:72:@41589.4]
  wire [7:0] _T_97298; // @[Mux.scala 19:72:@41596.4]
  wire [15:0] _T_97306; // @[Mux.scala 19:72:@41604.4]
  wire [15:0] _T_97308; // @[Mux.scala 19:72:@41605.4]
  wire [7:0] _T_97315; // @[Mux.scala 19:72:@41612.4]
  wire [15:0] _T_97323; // @[Mux.scala 19:72:@41620.4]
  wire [15:0] _T_97325; // @[Mux.scala 19:72:@41621.4]
  wire [7:0] _T_97332; // @[Mux.scala 19:72:@41628.4]
  wire [15:0] _T_97340; // @[Mux.scala 19:72:@41636.4]
  wire [15:0] _T_97342; // @[Mux.scala 19:72:@41637.4]
  wire [7:0] _T_97349; // @[Mux.scala 19:72:@41644.4]
  wire [15:0] _T_97357; // @[Mux.scala 19:72:@41652.4]
  wire [15:0] _T_97359; // @[Mux.scala 19:72:@41653.4]
  wire [7:0] _T_97366; // @[Mux.scala 19:72:@41660.4]
  wire [15:0] _T_97374; // @[Mux.scala 19:72:@41668.4]
  wire [15:0] _T_97376; // @[Mux.scala 19:72:@41669.4]
  wire [7:0] _T_97383; // @[Mux.scala 19:72:@41676.4]
  wire [15:0] _T_97391; // @[Mux.scala 19:72:@41684.4]
  wire [15:0] _T_97393; // @[Mux.scala 19:72:@41685.4]
  wire [7:0] _T_97400; // @[Mux.scala 19:72:@41692.4]
  wire [15:0] _T_97408; // @[Mux.scala 19:72:@41700.4]
  wire [15:0] _T_97410; // @[Mux.scala 19:72:@41701.4]
  wire [7:0] _T_97417; // @[Mux.scala 19:72:@41708.4]
  wire [15:0] _T_97425; // @[Mux.scala 19:72:@41716.4]
  wire [15:0] _T_97427; // @[Mux.scala 19:72:@41717.4]
  wire [7:0] _T_97434; // @[Mux.scala 19:72:@41724.4]
  wire [15:0] _T_97442; // @[Mux.scala 19:72:@41732.4]
  wire [15:0] _T_97444; // @[Mux.scala 19:72:@41733.4]
  wire [7:0] _T_97451; // @[Mux.scala 19:72:@41740.4]
  wire [15:0] _T_97459; // @[Mux.scala 19:72:@41748.4]
  wire [15:0] _T_97461; // @[Mux.scala 19:72:@41749.4]
  wire [7:0] _T_97468; // @[Mux.scala 19:72:@41756.4]
  wire [15:0] _T_97476; // @[Mux.scala 19:72:@41764.4]
  wire [15:0] _T_97478; // @[Mux.scala 19:72:@41765.4]
  wire [7:0] _T_97485; // @[Mux.scala 19:72:@41772.4]
  wire [15:0] _T_97493; // @[Mux.scala 19:72:@41780.4]
  wire [15:0] _T_97495; // @[Mux.scala 19:72:@41781.4]
  wire [7:0] _T_97502; // @[Mux.scala 19:72:@41788.4]
  wire [15:0] _T_97510; // @[Mux.scala 19:72:@41796.4]
  wire [15:0] _T_97512; // @[Mux.scala 19:72:@41797.4]
  wire [7:0] _T_97519; // @[Mux.scala 19:72:@41804.4]
  wire [15:0] _T_97527; // @[Mux.scala 19:72:@41812.4]
  wire [15:0] _T_97529; // @[Mux.scala 19:72:@41813.4]
  wire [7:0] _T_97536; // @[Mux.scala 19:72:@41820.4]
  wire [15:0] _T_97544; // @[Mux.scala 19:72:@41828.4]
  wire [15:0] _T_97546; // @[Mux.scala 19:72:@41829.4]
  wire [15:0] _T_97547; // @[Mux.scala 19:72:@41830.4]
  wire [15:0] _T_97548; // @[Mux.scala 19:72:@41831.4]
  wire [15:0] _T_97549; // @[Mux.scala 19:72:@41832.4]
  wire [15:0] _T_97550; // @[Mux.scala 19:72:@41833.4]
  wire [15:0] _T_97551; // @[Mux.scala 19:72:@41834.4]
  wire [15:0] _T_97552; // @[Mux.scala 19:72:@41835.4]
  wire [15:0] _T_97553; // @[Mux.scala 19:72:@41836.4]
  wire [15:0] _T_97554; // @[Mux.scala 19:72:@41837.4]
  wire [15:0] _T_97555; // @[Mux.scala 19:72:@41838.4]
  wire [15:0] _T_97556; // @[Mux.scala 19:72:@41839.4]
  wire [15:0] _T_97557; // @[Mux.scala 19:72:@41840.4]
  wire [15:0] _T_97558; // @[Mux.scala 19:72:@41841.4]
  wire [15:0] _T_97559; // @[Mux.scala 19:72:@41842.4]
  wire [15:0] _T_97560; // @[Mux.scala 19:72:@41843.4]
  wire [15:0] _T_97561; // @[Mux.scala 19:72:@41844.4]
  wire  outputPriorityPorts_0_0; // @[Mux.scala 19:72:@41848.4]
  wire  outputPriorityPorts_0_1; // @[Mux.scala 19:72:@41850.4]
  wire  outputPriorityPorts_0_2; // @[Mux.scala 19:72:@41852.4]
  wire  outputPriorityPorts_0_3; // @[Mux.scala 19:72:@41854.4]
  wire  outputPriorityPorts_0_4; // @[Mux.scala 19:72:@41856.4]
  wire  outputPriorityPorts_0_5; // @[Mux.scala 19:72:@41858.4]
  wire  outputPriorityPorts_0_6; // @[Mux.scala 19:72:@41860.4]
  wire  outputPriorityPorts_0_7; // @[Mux.scala 19:72:@41862.4]
  wire  outputPriorityPorts_0_8; // @[Mux.scala 19:72:@41864.4]
  wire  outputPriorityPorts_0_9; // @[Mux.scala 19:72:@41866.4]
  wire  outputPriorityPorts_0_10; // @[Mux.scala 19:72:@41868.4]
  wire  outputPriorityPorts_0_11; // @[Mux.scala 19:72:@41870.4]
  wire  outputPriorityPorts_0_12; // @[Mux.scala 19:72:@41872.4]
  wire  outputPriorityPorts_0_13; // @[Mux.scala 19:72:@41874.4]
  wire  outputPriorityPorts_0_14; // @[Mux.scala 19:72:@41876.4]
  wire  outputPriorityPorts_0_15; // @[Mux.scala 19:72:@41878.4]
  wire  _T_97704; // @[AxiLoadQueue.scala 315:47:@41900.6]
  wire [30:0] _GEN_2128; // @[AxiLoadQueue.scala 316:36:@41904.6]
  wire  _GEN_2129; // @[AxiLoadQueue.scala 316:36:@41904.6]
  wire  _GEN_2130; // @[AxiLoadQueue.scala 310:34:@41896.4]
  wire [30:0] _GEN_2131; // @[AxiLoadQueue.scala 310:34:@41896.4]
  wire  _T_97719; // @[AxiLoadQueue.scala 315:47:@41913.6]
  wire [30:0] _GEN_2132; // @[AxiLoadQueue.scala 316:36:@41917.6]
  wire  _GEN_2133; // @[AxiLoadQueue.scala 316:36:@41917.6]
  wire  _GEN_2134; // @[AxiLoadQueue.scala 310:34:@41909.4]
  wire [30:0] _GEN_2135; // @[AxiLoadQueue.scala 310:34:@41909.4]
  wire  _T_97734; // @[AxiLoadQueue.scala 315:47:@41926.6]
  wire [30:0] _GEN_2136; // @[AxiLoadQueue.scala 316:36:@41930.6]
  wire  _GEN_2137; // @[AxiLoadQueue.scala 316:36:@41930.6]
  wire  _GEN_2138; // @[AxiLoadQueue.scala 310:34:@41922.4]
  wire [30:0] _GEN_2139; // @[AxiLoadQueue.scala 310:34:@41922.4]
  wire  _T_97749; // @[AxiLoadQueue.scala 315:47:@41939.6]
  wire [30:0] _GEN_2140; // @[AxiLoadQueue.scala 316:36:@41943.6]
  wire  _GEN_2141; // @[AxiLoadQueue.scala 316:36:@41943.6]
  wire  _GEN_2142; // @[AxiLoadQueue.scala 310:34:@41935.4]
  wire [30:0] _GEN_2143; // @[AxiLoadQueue.scala 310:34:@41935.4]
  wire  _T_97764; // @[AxiLoadQueue.scala 315:47:@41952.6]
  wire [30:0] _GEN_2144; // @[AxiLoadQueue.scala 316:36:@41956.6]
  wire  _GEN_2145; // @[AxiLoadQueue.scala 316:36:@41956.6]
  wire  _GEN_2146; // @[AxiLoadQueue.scala 310:34:@41948.4]
  wire [30:0] _GEN_2147; // @[AxiLoadQueue.scala 310:34:@41948.4]
  wire  _T_97779; // @[AxiLoadQueue.scala 315:47:@41965.6]
  wire [30:0] _GEN_2148; // @[AxiLoadQueue.scala 316:36:@41969.6]
  wire  _GEN_2149; // @[AxiLoadQueue.scala 316:36:@41969.6]
  wire  _GEN_2150; // @[AxiLoadQueue.scala 310:34:@41961.4]
  wire [30:0] _GEN_2151; // @[AxiLoadQueue.scala 310:34:@41961.4]
  wire  _T_97794; // @[AxiLoadQueue.scala 315:47:@41978.6]
  wire [30:0] _GEN_2152; // @[AxiLoadQueue.scala 316:36:@41982.6]
  wire  _GEN_2153; // @[AxiLoadQueue.scala 316:36:@41982.6]
  wire  _GEN_2154; // @[AxiLoadQueue.scala 310:34:@41974.4]
  wire [30:0] _GEN_2155; // @[AxiLoadQueue.scala 310:34:@41974.4]
  wire  _T_97809; // @[AxiLoadQueue.scala 315:47:@41991.6]
  wire [30:0] _GEN_2156; // @[AxiLoadQueue.scala 316:36:@41995.6]
  wire  _GEN_2157; // @[AxiLoadQueue.scala 316:36:@41995.6]
  wire  _GEN_2158; // @[AxiLoadQueue.scala 310:34:@41987.4]
  wire [30:0] _GEN_2159; // @[AxiLoadQueue.scala 310:34:@41987.4]
  wire  _T_97824; // @[AxiLoadQueue.scala 315:47:@42004.6]
  wire [30:0] _GEN_2160; // @[AxiLoadQueue.scala 316:36:@42008.6]
  wire  _GEN_2161; // @[AxiLoadQueue.scala 316:36:@42008.6]
  wire  _GEN_2162; // @[AxiLoadQueue.scala 310:34:@42000.4]
  wire [30:0] _GEN_2163; // @[AxiLoadQueue.scala 310:34:@42000.4]
  wire  _T_97839; // @[AxiLoadQueue.scala 315:47:@42017.6]
  wire [30:0] _GEN_2164; // @[AxiLoadQueue.scala 316:36:@42021.6]
  wire  _GEN_2165; // @[AxiLoadQueue.scala 316:36:@42021.6]
  wire  _GEN_2166; // @[AxiLoadQueue.scala 310:34:@42013.4]
  wire [30:0] _GEN_2167; // @[AxiLoadQueue.scala 310:34:@42013.4]
  wire  _T_97854; // @[AxiLoadQueue.scala 315:47:@42030.6]
  wire [30:0] _GEN_2168; // @[AxiLoadQueue.scala 316:36:@42034.6]
  wire  _GEN_2169; // @[AxiLoadQueue.scala 316:36:@42034.6]
  wire  _GEN_2170; // @[AxiLoadQueue.scala 310:34:@42026.4]
  wire [30:0] _GEN_2171; // @[AxiLoadQueue.scala 310:34:@42026.4]
  wire  _T_97869; // @[AxiLoadQueue.scala 315:47:@42043.6]
  wire [30:0] _GEN_2172; // @[AxiLoadQueue.scala 316:36:@42047.6]
  wire  _GEN_2173; // @[AxiLoadQueue.scala 316:36:@42047.6]
  wire  _GEN_2174; // @[AxiLoadQueue.scala 310:34:@42039.4]
  wire [30:0] _GEN_2175; // @[AxiLoadQueue.scala 310:34:@42039.4]
  wire  _T_97884; // @[AxiLoadQueue.scala 315:47:@42056.6]
  wire [30:0] _GEN_2176; // @[AxiLoadQueue.scala 316:36:@42060.6]
  wire  _GEN_2177; // @[AxiLoadQueue.scala 316:36:@42060.6]
  wire  _GEN_2178; // @[AxiLoadQueue.scala 310:34:@42052.4]
  wire [30:0] _GEN_2179; // @[AxiLoadQueue.scala 310:34:@42052.4]
  wire  _T_97899; // @[AxiLoadQueue.scala 315:47:@42069.6]
  wire [30:0] _GEN_2180; // @[AxiLoadQueue.scala 316:36:@42073.6]
  wire  _GEN_2181; // @[AxiLoadQueue.scala 316:36:@42073.6]
  wire  _GEN_2182; // @[AxiLoadQueue.scala 310:34:@42065.4]
  wire [30:0] _GEN_2183; // @[AxiLoadQueue.scala 310:34:@42065.4]
  wire  _T_97914; // @[AxiLoadQueue.scala 315:47:@42082.6]
  wire [30:0] _GEN_2184; // @[AxiLoadQueue.scala 316:36:@42086.6]
  wire  _GEN_2185; // @[AxiLoadQueue.scala 316:36:@42086.6]
  wire  _GEN_2186; // @[AxiLoadQueue.scala 310:34:@42078.4]
  wire [30:0] _GEN_2187; // @[AxiLoadQueue.scala 310:34:@42078.4]
  wire  _T_97929; // @[AxiLoadQueue.scala 315:47:@42095.6]
  wire [30:0] _GEN_2188; // @[AxiLoadQueue.scala 316:36:@42099.6]
  wire  _GEN_2189; // @[AxiLoadQueue.scala 316:36:@42099.6]
  wire  _GEN_2190; // @[AxiLoadQueue.scala 310:34:@42091.4]
  wire [30:0] _GEN_2191; // @[AxiLoadQueue.scala 310:34:@42091.4]
  wire  _T_97964; // @[AxiLoadQueue.scala 328:108:@42105.4]
  wire  _T_97966; // @[AxiLoadQueue.scala 329:34:@42106.4]
  wire  _T_97967; // @[AxiLoadQueue.scala 329:31:@42107.4]
  wire  loadCompleting_0; // @[AxiLoadQueue.scala 329:63:@42108.4]
  wire  _T_97978; // @[AxiLoadQueue.scala 328:108:@42113.4]
  wire  _T_97980; // @[AxiLoadQueue.scala 329:34:@42114.4]
  wire  _T_97981; // @[AxiLoadQueue.scala 329:31:@42115.4]
  wire  loadCompleting_1; // @[AxiLoadQueue.scala 329:63:@42116.4]
  wire  _T_97992; // @[AxiLoadQueue.scala 328:108:@42121.4]
  wire  _T_97994; // @[AxiLoadQueue.scala 329:34:@42122.4]
  wire  _T_97995; // @[AxiLoadQueue.scala 329:31:@42123.4]
  wire  loadCompleting_2; // @[AxiLoadQueue.scala 329:63:@42124.4]
  wire  _T_98006; // @[AxiLoadQueue.scala 328:108:@42129.4]
  wire  _T_98008; // @[AxiLoadQueue.scala 329:34:@42130.4]
  wire  _T_98009; // @[AxiLoadQueue.scala 329:31:@42131.4]
  wire  loadCompleting_3; // @[AxiLoadQueue.scala 329:63:@42132.4]
  wire  _T_98020; // @[AxiLoadQueue.scala 328:108:@42137.4]
  wire  _T_98022; // @[AxiLoadQueue.scala 329:34:@42138.4]
  wire  _T_98023; // @[AxiLoadQueue.scala 329:31:@42139.4]
  wire  loadCompleting_4; // @[AxiLoadQueue.scala 329:63:@42140.4]
  wire  _T_98034; // @[AxiLoadQueue.scala 328:108:@42145.4]
  wire  _T_98036; // @[AxiLoadQueue.scala 329:34:@42146.4]
  wire  _T_98037; // @[AxiLoadQueue.scala 329:31:@42147.4]
  wire  loadCompleting_5; // @[AxiLoadQueue.scala 329:63:@42148.4]
  wire  _T_98048; // @[AxiLoadQueue.scala 328:108:@42153.4]
  wire  _T_98050; // @[AxiLoadQueue.scala 329:34:@42154.4]
  wire  _T_98051; // @[AxiLoadQueue.scala 329:31:@42155.4]
  wire  loadCompleting_6; // @[AxiLoadQueue.scala 329:63:@42156.4]
  wire  _T_98062; // @[AxiLoadQueue.scala 328:108:@42161.4]
  wire  _T_98064; // @[AxiLoadQueue.scala 329:34:@42162.4]
  wire  _T_98065; // @[AxiLoadQueue.scala 329:31:@42163.4]
  wire  loadCompleting_7; // @[AxiLoadQueue.scala 329:63:@42164.4]
  wire  _T_98076; // @[AxiLoadQueue.scala 328:108:@42169.4]
  wire  _T_98078; // @[AxiLoadQueue.scala 329:34:@42170.4]
  wire  _T_98079; // @[AxiLoadQueue.scala 329:31:@42171.4]
  wire  loadCompleting_8; // @[AxiLoadQueue.scala 329:63:@42172.4]
  wire  _T_98090; // @[AxiLoadQueue.scala 328:108:@42177.4]
  wire  _T_98092; // @[AxiLoadQueue.scala 329:34:@42178.4]
  wire  _T_98093; // @[AxiLoadQueue.scala 329:31:@42179.4]
  wire  loadCompleting_9; // @[AxiLoadQueue.scala 329:63:@42180.4]
  wire  _T_98104; // @[AxiLoadQueue.scala 328:108:@42185.4]
  wire  _T_98106; // @[AxiLoadQueue.scala 329:34:@42186.4]
  wire  _T_98107; // @[AxiLoadQueue.scala 329:31:@42187.4]
  wire  loadCompleting_10; // @[AxiLoadQueue.scala 329:63:@42188.4]
  wire  _T_98118; // @[AxiLoadQueue.scala 328:108:@42193.4]
  wire  _T_98120; // @[AxiLoadQueue.scala 329:34:@42194.4]
  wire  _T_98121; // @[AxiLoadQueue.scala 329:31:@42195.4]
  wire  loadCompleting_11; // @[AxiLoadQueue.scala 329:63:@42196.4]
  wire  _T_98132; // @[AxiLoadQueue.scala 328:108:@42201.4]
  wire  _T_98134; // @[AxiLoadQueue.scala 329:34:@42202.4]
  wire  _T_98135; // @[AxiLoadQueue.scala 329:31:@42203.4]
  wire  loadCompleting_12; // @[AxiLoadQueue.scala 329:63:@42204.4]
  wire  _T_98146; // @[AxiLoadQueue.scala 328:108:@42209.4]
  wire  _T_98148; // @[AxiLoadQueue.scala 329:34:@42210.4]
  wire  _T_98149; // @[AxiLoadQueue.scala 329:31:@42211.4]
  wire  loadCompleting_13; // @[AxiLoadQueue.scala 329:63:@42212.4]
  wire  _T_98160; // @[AxiLoadQueue.scala 328:108:@42217.4]
  wire  _T_98162; // @[AxiLoadQueue.scala 329:34:@42218.4]
  wire  _T_98163; // @[AxiLoadQueue.scala 329:31:@42219.4]
  wire  loadCompleting_14; // @[AxiLoadQueue.scala 329:63:@42220.4]
  wire  _T_98174; // @[AxiLoadQueue.scala 328:108:@42225.4]
  wire  _T_98176; // @[AxiLoadQueue.scala 329:34:@42226.4]
  wire  _T_98177; // @[AxiLoadQueue.scala 329:31:@42227.4]
  wire  loadCompleting_15; // @[AxiLoadQueue.scala 329:63:@42228.4]
  wire  _GEN_2192; // @[AxiLoadQueue.scala 339:46:@42237.6]
  wire  _GEN_2193; // @[AxiLoadQueue.scala 337:34:@42233.4]
  wire  _GEN_2194; // @[AxiLoadQueue.scala 339:46:@42244.6]
  wire  _GEN_2195; // @[AxiLoadQueue.scala 337:34:@42240.4]
  wire  _GEN_2196; // @[AxiLoadQueue.scala 339:46:@42251.6]
  wire  _GEN_2197; // @[AxiLoadQueue.scala 337:34:@42247.4]
  wire  _GEN_2198; // @[AxiLoadQueue.scala 339:46:@42258.6]
  wire  _GEN_2199; // @[AxiLoadQueue.scala 337:34:@42254.4]
  wire  _GEN_2200; // @[AxiLoadQueue.scala 339:46:@42265.6]
  wire  _GEN_2201; // @[AxiLoadQueue.scala 337:34:@42261.4]
  wire  _GEN_2202; // @[AxiLoadQueue.scala 339:46:@42272.6]
  wire  _GEN_2203; // @[AxiLoadQueue.scala 337:34:@42268.4]
  wire  _GEN_2204; // @[AxiLoadQueue.scala 339:46:@42279.6]
  wire  _GEN_2205; // @[AxiLoadQueue.scala 337:34:@42275.4]
  wire  _GEN_2206; // @[AxiLoadQueue.scala 339:46:@42286.6]
  wire  _GEN_2207; // @[AxiLoadQueue.scala 337:34:@42282.4]
  wire  _GEN_2208; // @[AxiLoadQueue.scala 339:46:@42293.6]
  wire  _GEN_2209; // @[AxiLoadQueue.scala 337:34:@42289.4]
  wire  _GEN_2210; // @[AxiLoadQueue.scala 339:46:@42300.6]
  wire  _GEN_2211; // @[AxiLoadQueue.scala 337:34:@42296.4]
  wire  _GEN_2212; // @[AxiLoadQueue.scala 339:46:@42307.6]
  wire  _GEN_2213; // @[AxiLoadQueue.scala 337:34:@42303.4]
  wire  _GEN_2214; // @[AxiLoadQueue.scala 339:46:@42314.6]
  wire  _GEN_2215; // @[AxiLoadQueue.scala 337:34:@42310.4]
  wire  _GEN_2216; // @[AxiLoadQueue.scala 339:46:@42321.6]
  wire  _GEN_2217; // @[AxiLoadQueue.scala 337:34:@42317.4]
  wire  _GEN_2218; // @[AxiLoadQueue.scala 339:46:@42328.6]
  wire  _GEN_2219; // @[AxiLoadQueue.scala 337:34:@42324.4]
  wire  _GEN_2220; // @[AxiLoadQueue.scala 339:46:@42335.6]
  wire  _GEN_2221; // @[AxiLoadQueue.scala 337:34:@42331.4]
  wire  _GEN_2222; // @[AxiLoadQueue.scala 339:46:@42342.6]
  wire  _GEN_2223; // @[AxiLoadQueue.scala 337:34:@42338.4]
  wire  _T_98308; // @[AxiLoadQueue.scala 350:24:@42411.4]
  wire  _T_98309; // @[AxiLoadQueue.scala 350:24:@42412.4]
  wire  _T_98310; // @[AxiLoadQueue.scala 350:24:@42413.4]
  wire  _T_98311; // @[AxiLoadQueue.scala 350:24:@42414.4]
  wire  _T_98312; // @[AxiLoadQueue.scala 350:24:@42415.4]
  wire  _T_98313; // @[AxiLoadQueue.scala 350:24:@42416.4]
  wire  _T_98314; // @[AxiLoadQueue.scala 350:24:@42417.4]
  wire  _T_98315; // @[AxiLoadQueue.scala 350:24:@42418.4]
  wire  _T_98316; // @[AxiLoadQueue.scala 350:24:@42419.4]
  wire  _T_98317; // @[AxiLoadQueue.scala 350:24:@42420.4]
  wire  _T_98318; // @[AxiLoadQueue.scala 350:24:@42421.4]
  wire  _T_98319; // @[AxiLoadQueue.scala 350:24:@42422.4]
  wire  _T_98320; // @[AxiLoadQueue.scala 350:24:@42423.4]
  wire  _T_98321; // @[AxiLoadQueue.scala 350:24:@42424.4]
  wire  _T_98322; // @[AxiLoadQueue.scala 350:24:@42425.4]
  wire [3:0] _T_98339; // @[Mux.scala 31:69:@42427.6]
  wire [3:0] _T_98340; // @[Mux.scala 31:69:@42428.6]
  wire [3:0] _T_98341; // @[Mux.scala 31:69:@42429.6]
  wire [3:0] _T_98342; // @[Mux.scala 31:69:@42430.6]
  wire [3:0] _T_98343; // @[Mux.scala 31:69:@42431.6]
  wire [3:0] _T_98344; // @[Mux.scala 31:69:@42432.6]
  wire [3:0] _T_98345; // @[Mux.scala 31:69:@42433.6]
  wire [3:0] _T_98346; // @[Mux.scala 31:69:@42434.6]
  wire [3:0] _T_98347; // @[Mux.scala 31:69:@42435.6]
  wire [3:0] _T_98348; // @[Mux.scala 31:69:@42436.6]
  wire [3:0] _T_98349; // @[Mux.scala 31:69:@42437.6]
  wire [3:0] _T_98350; // @[Mux.scala 31:69:@42438.6]
  wire [3:0] _T_98351; // @[Mux.scala 31:69:@42439.6]
  wire [3:0] _T_98352; // @[Mux.scala 31:69:@42440.6]
  wire [3:0] _T_98353; // @[Mux.scala 31:69:@42441.6]
  wire [31:0] _GEN_2225; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2226; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2227; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2228; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2229; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2230; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2231; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2232; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2233; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2234; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2235; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2236; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2237; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2238; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire [31:0] _GEN_2239; // @[AxiLoadQueue.scala 351:37:@42442.6]
  wire  _GEN_2243; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2244; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2245; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2246; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2247; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2248; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2249; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2250; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2251; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2252; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2253; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2254; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2255; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2256; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2257; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2259; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2260; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2261; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2262; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2263; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2264; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2265; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2266; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2267; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2268; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2269; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2270; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2271; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2272; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _GEN_2273; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _T_98364; // @[AxiLoadQueue.scala 365:29:@42449.4]
  wire  _T_98365; // @[AxiLoadQueue.scala 365:63:@42450.4]
  wire  _T_98367; // @[AxiLoadQueue.scala 365:75:@42451.4]
  wire  _T_98368; // @[AxiLoadQueue.scala 365:72:@42452.4]
  wire  _T_98369; // @[AxiLoadQueue.scala 365:54:@42453.4]
  wire [4:0] _T_98372; // @[util.scala 10:8:@42455.6]
  wire [4:0] _GEN_64; // @[util.scala 10:14:@42456.6]
  wire [4:0] _T_98373; // @[util.scala 10:14:@42456.6]
  wire [4:0] _GEN_2274; // @[AxiLoadQueue.scala 365:91:@42454.4]
  wire [3:0] _GEN_2372; // @[util.scala 10:8:@42460.6]
  wire [4:0] _T_98375; // @[util.scala 10:8:@42460.6]
  wire [4:0] _GEN_65; // @[util.scala 10:14:@42461.6]
  wire [4:0] _T_98376; // @[util.scala 10:14:@42461.6]
  wire [4:0] _GEN_2275; // @[AxiLoadQueue.scala 369:20:@42459.4]
  wire  _T_98378; // @[AxiLoadQueue.scala 373:82:@42464.4]
  wire  _T_98379; // @[AxiLoadQueue.scala 373:79:@42465.4]
  wire  _T_98381; // @[AxiLoadQueue.scala 373:82:@42466.4]
  wire  _T_98382; // @[AxiLoadQueue.scala 373:79:@42467.4]
  wire  _T_98384; // @[AxiLoadQueue.scala 373:82:@42468.4]
  wire  _T_98385; // @[AxiLoadQueue.scala 373:79:@42469.4]
  wire  _T_98387; // @[AxiLoadQueue.scala 373:82:@42470.4]
  wire  _T_98388; // @[AxiLoadQueue.scala 373:79:@42471.4]
  wire  _T_98390; // @[AxiLoadQueue.scala 373:82:@42472.4]
  wire  _T_98391; // @[AxiLoadQueue.scala 373:79:@42473.4]
  wire  _T_98393; // @[AxiLoadQueue.scala 373:82:@42474.4]
  wire  _T_98394; // @[AxiLoadQueue.scala 373:79:@42475.4]
  wire  _T_98396; // @[AxiLoadQueue.scala 373:82:@42476.4]
  wire  _T_98397; // @[AxiLoadQueue.scala 373:79:@42477.4]
  wire  _T_98399; // @[AxiLoadQueue.scala 373:82:@42478.4]
  wire  _T_98400; // @[AxiLoadQueue.scala 373:79:@42479.4]
  wire  _T_98402; // @[AxiLoadQueue.scala 373:82:@42480.4]
  wire  _T_98403; // @[AxiLoadQueue.scala 373:79:@42481.4]
  wire  _T_98405; // @[AxiLoadQueue.scala 373:82:@42482.4]
  wire  _T_98406; // @[AxiLoadQueue.scala 373:79:@42483.4]
  wire  _T_98408; // @[AxiLoadQueue.scala 373:82:@42484.4]
  wire  _T_98409; // @[AxiLoadQueue.scala 373:79:@42485.4]
  wire  _T_98411; // @[AxiLoadQueue.scala 373:82:@42486.4]
  wire  _T_98412; // @[AxiLoadQueue.scala 373:79:@42487.4]
  wire  _T_98414; // @[AxiLoadQueue.scala 373:82:@42488.4]
  wire  _T_98415; // @[AxiLoadQueue.scala 373:79:@42489.4]
  wire  _T_98417; // @[AxiLoadQueue.scala 373:82:@42490.4]
  wire  _T_98418; // @[AxiLoadQueue.scala 373:79:@42491.4]
  wire  _T_98420; // @[AxiLoadQueue.scala 373:82:@42492.4]
  wire  _T_98421; // @[AxiLoadQueue.scala 373:79:@42493.4]
  wire  _T_98423; // @[AxiLoadQueue.scala 373:82:@42494.4]
  wire  _T_98424; // @[AxiLoadQueue.scala 373:79:@42495.4]
  wire  _T_98449; // @[AxiLoadQueue.scala 373:96:@42514.4]
  wire  _T_98450; // @[AxiLoadQueue.scala 373:96:@42515.4]
  wire  _T_98451; // @[AxiLoadQueue.scala 373:96:@42516.4]
  wire  _T_98452; // @[AxiLoadQueue.scala 373:96:@42517.4]
  wire  _T_98453; // @[AxiLoadQueue.scala 373:96:@42518.4]
  wire  _T_98454; // @[AxiLoadQueue.scala 373:96:@42519.4]
  wire  _T_98455; // @[AxiLoadQueue.scala 373:96:@42520.4]
  wire  _T_98456; // @[AxiLoadQueue.scala 373:96:@42521.4]
  wire  _T_98457; // @[AxiLoadQueue.scala 373:96:@42522.4]
  wire  _T_98458; // @[AxiLoadQueue.scala 373:96:@42523.4]
  wire  _T_98459; // @[AxiLoadQueue.scala 373:96:@42524.4]
  wire  _T_98460; // @[AxiLoadQueue.scala 373:96:@42525.4]
  wire  _T_98461; // @[AxiLoadQueue.scala 373:96:@42526.4]
  wire  _T_98462; // @[AxiLoadQueue.scala 373:96:@42527.4]
  assign _GEN_2276 = {{2'd0}, tail}; // @[util.scala 14:20:@5026.4]
  assign _T_1722 = 6'h10 - _GEN_2276; // @[util.scala 14:20:@5026.4]
  assign _T_1723 = $unsigned(_T_1722); // @[util.scala 14:20:@5027.4]
  assign _T_1724 = _T_1723[5:0]; // @[util.scala 14:20:@5028.4]
  assign _GEN_0 = _T_1724 % 6'h10; // @[util.scala 14:25:@5029.4]
  assign _T_1725 = _GEN_0[4:0]; // @[util.scala 14:25:@5029.4]
  assign _GEN_2277 = {{4'd0}, io_bbNumLoads}; // @[AxiLoadQueue.scala 71:46:@5030.4]
  assign _T_1726 = _T_1725 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5030.4]
  assign initBits_0 = _T_1726 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5031.4]
  assign _T_1731 = 6'h11 - _GEN_2276; // @[util.scala 14:20:@5033.4]
  assign _T_1732 = $unsigned(_T_1731); // @[util.scala 14:20:@5034.4]
  assign _T_1733 = _T_1732[5:0]; // @[util.scala 14:20:@5035.4]
  assign _GEN_16 = _T_1733 % 6'h10; // @[util.scala 14:25:@5036.4]
  assign _T_1734 = _GEN_16[4:0]; // @[util.scala 14:25:@5036.4]
  assign _T_1735 = _T_1734 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5037.4]
  assign initBits_1 = _T_1735 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5038.4]
  assign _T_1740 = 6'h12 - _GEN_2276; // @[util.scala 14:20:@5040.4]
  assign _T_1741 = $unsigned(_T_1740); // @[util.scala 14:20:@5041.4]
  assign _T_1742 = _T_1741[5:0]; // @[util.scala 14:20:@5042.4]
  assign _GEN_17 = _T_1742 % 6'h10; // @[util.scala 14:25:@5043.4]
  assign _T_1743 = _GEN_17[4:0]; // @[util.scala 14:25:@5043.4]
  assign _T_1744 = _T_1743 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5044.4]
  assign initBits_2 = _T_1744 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5045.4]
  assign _T_1749 = 6'h13 - _GEN_2276; // @[util.scala 14:20:@5047.4]
  assign _T_1750 = $unsigned(_T_1749); // @[util.scala 14:20:@5048.4]
  assign _T_1751 = _T_1750[5:0]; // @[util.scala 14:20:@5049.4]
  assign _GEN_18 = _T_1751 % 6'h10; // @[util.scala 14:25:@5050.4]
  assign _T_1752 = _GEN_18[4:0]; // @[util.scala 14:25:@5050.4]
  assign _T_1753 = _T_1752 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5051.4]
  assign initBits_3 = _T_1753 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5052.4]
  assign _T_1758 = 6'h14 - _GEN_2276; // @[util.scala 14:20:@5054.4]
  assign _T_1759 = $unsigned(_T_1758); // @[util.scala 14:20:@5055.4]
  assign _T_1760 = _T_1759[5:0]; // @[util.scala 14:20:@5056.4]
  assign _GEN_19 = _T_1760 % 6'h10; // @[util.scala 14:25:@5057.4]
  assign _T_1761 = _GEN_19[4:0]; // @[util.scala 14:25:@5057.4]
  assign _T_1762 = _T_1761 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5058.4]
  assign initBits_4 = _T_1762 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5059.4]
  assign _T_1767 = 6'h15 - _GEN_2276; // @[util.scala 14:20:@5061.4]
  assign _T_1768 = $unsigned(_T_1767); // @[util.scala 14:20:@5062.4]
  assign _T_1769 = _T_1768[5:0]; // @[util.scala 14:20:@5063.4]
  assign _GEN_20 = _T_1769 % 6'h10; // @[util.scala 14:25:@5064.4]
  assign _T_1770 = _GEN_20[4:0]; // @[util.scala 14:25:@5064.4]
  assign _T_1771 = _T_1770 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5065.4]
  assign initBits_5 = _T_1771 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5066.4]
  assign _T_1776 = 6'h16 - _GEN_2276; // @[util.scala 14:20:@5068.4]
  assign _T_1777 = $unsigned(_T_1776); // @[util.scala 14:20:@5069.4]
  assign _T_1778 = _T_1777[5:0]; // @[util.scala 14:20:@5070.4]
  assign _GEN_21 = _T_1778 % 6'h10; // @[util.scala 14:25:@5071.4]
  assign _T_1779 = _GEN_21[4:0]; // @[util.scala 14:25:@5071.4]
  assign _T_1780 = _T_1779 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5072.4]
  assign initBits_6 = _T_1780 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5073.4]
  assign _T_1785 = 6'h17 - _GEN_2276; // @[util.scala 14:20:@5075.4]
  assign _T_1786 = $unsigned(_T_1785); // @[util.scala 14:20:@5076.4]
  assign _T_1787 = _T_1786[5:0]; // @[util.scala 14:20:@5077.4]
  assign _GEN_22 = _T_1787 % 6'h10; // @[util.scala 14:25:@5078.4]
  assign _T_1788 = _GEN_22[4:0]; // @[util.scala 14:25:@5078.4]
  assign _T_1789 = _T_1788 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5079.4]
  assign initBits_7 = _T_1789 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5080.4]
  assign _T_1794 = 6'h18 - _GEN_2276; // @[util.scala 14:20:@5082.4]
  assign _T_1795 = $unsigned(_T_1794); // @[util.scala 14:20:@5083.4]
  assign _T_1796 = _T_1795[5:0]; // @[util.scala 14:20:@5084.4]
  assign _GEN_23 = _T_1796 % 6'h10; // @[util.scala 14:25:@5085.4]
  assign _T_1797 = _GEN_23[4:0]; // @[util.scala 14:25:@5085.4]
  assign _T_1798 = _T_1797 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5086.4]
  assign initBits_8 = _T_1798 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5087.4]
  assign _T_1803 = 6'h19 - _GEN_2276; // @[util.scala 14:20:@5089.4]
  assign _T_1804 = $unsigned(_T_1803); // @[util.scala 14:20:@5090.4]
  assign _T_1805 = _T_1804[5:0]; // @[util.scala 14:20:@5091.4]
  assign _GEN_24 = _T_1805 % 6'h10; // @[util.scala 14:25:@5092.4]
  assign _T_1806 = _GEN_24[4:0]; // @[util.scala 14:25:@5092.4]
  assign _T_1807 = _T_1806 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5093.4]
  assign initBits_9 = _T_1807 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5094.4]
  assign _T_1812 = 6'h1a - _GEN_2276; // @[util.scala 14:20:@5096.4]
  assign _T_1813 = $unsigned(_T_1812); // @[util.scala 14:20:@5097.4]
  assign _T_1814 = _T_1813[5:0]; // @[util.scala 14:20:@5098.4]
  assign _GEN_25 = _T_1814 % 6'h10; // @[util.scala 14:25:@5099.4]
  assign _T_1815 = _GEN_25[4:0]; // @[util.scala 14:25:@5099.4]
  assign _T_1816 = _T_1815 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5100.4]
  assign initBits_10 = _T_1816 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5101.4]
  assign _T_1821 = 6'h1b - _GEN_2276; // @[util.scala 14:20:@5103.4]
  assign _T_1822 = $unsigned(_T_1821); // @[util.scala 14:20:@5104.4]
  assign _T_1823 = _T_1822[5:0]; // @[util.scala 14:20:@5105.4]
  assign _GEN_26 = _T_1823 % 6'h10; // @[util.scala 14:25:@5106.4]
  assign _T_1824 = _GEN_26[4:0]; // @[util.scala 14:25:@5106.4]
  assign _T_1825 = _T_1824 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5107.4]
  assign initBits_11 = _T_1825 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5108.4]
  assign _T_1830 = 6'h1c - _GEN_2276; // @[util.scala 14:20:@5110.4]
  assign _T_1831 = $unsigned(_T_1830); // @[util.scala 14:20:@5111.4]
  assign _T_1832 = _T_1831[5:0]; // @[util.scala 14:20:@5112.4]
  assign _GEN_27 = _T_1832 % 6'h10; // @[util.scala 14:25:@5113.4]
  assign _T_1833 = _GEN_27[4:0]; // @[util.scala 14:25:@5113.4]
  assign _T_1834 = _T_1833 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5114.4]
  assign initBits_12 = _T_1834 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5115.4]
  assign _T_1839 = 6'h1d - _GEN_2276; // @[util.scala 14:20:@5117.4]
  assign _T_1840 = $unsigned(_T_1839); // @[util.scala 14:20:@5118.4]
  assign _T_1841 = _T_1840[5:0]; // @[util.scala 14:20:@5119.4]
  assign _GEN_28 = _T_1841 % 6'h10; // @[util.scala 14:25:@5120.4]
  assign _T_1842 = _GEN_28[4:0]; // @[util.scala 14:25:@5120.4]
  assign _T_1843 = _T_1842 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5121.4]
  assign initBits_13 = _T_1843 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5122.4]
  assign _T_1848 = 6'h1e - _GEN_2276; // @[util.scala 14:20:@5124.4]
  assign _T_1849 = $unsigned(_T_1848); // @[util.scala 14:20:@5125.4]
  assign _T_1850 = _T_1849[5:0]; // @[util.scala 14:20:@5126.4]
  assign _GEN_29 = _T_1850 % 6'h10; // @[util.scala 14:25:@5127.4]
  assign _T_1851 = _GEN_29[4:0]; // @[util.scala 14:25:@5127.4]
  assign _T_1852 = _T_1851 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5128.4]
  assign initBits_14 = _T_1852 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5129.4]
  assign _T_1857 = 6'h1f - _GEN_2276; // @[util.scala 14:20:@5131.4]
  assign _T_1858 = $unsigned(_T_1857); // @[util.scala 14:20:@5132.4]
  assign _T_1859 = _T_1858[5:0]; // @[util.scala 14:20:@5133.4]
  assign _GEN_30 = _T_1859 % 6'h10; // @[util.scala 14:25:@5134.4]
  assign _T_1860 = _GEN_30[4:0]; // @[util.scala 14:25:@5134.4]
  assign _T_1861 = _T_1860 < _GEN_2277; // @[AxiLoadQueue.scala 71:46:@5135.4]
  assign initBits_15 = _T_1861 & io_bbStart; // @[AxiLoadQueue.scala 71:63:@5136.4]
  assign _T_1884 = allocatedEntries_0 | initBits_0; // @[AxiLoadQueue.scala 73:78:@5154.4]
  assign _T_1885 = allocatedEntries_1 | initBits_1; // @[AxiLoadQueue.scala 73:78:@5155.4]
  assign _T_1886 = allocatedEntries_2 | initBits_2; // @[AxiLoadQueue.scala 73:78:@5156.4]
  assign _T_1887 = allocatedEntries_3 | initBits_3; // @[AxiLoadQueue.scala 73:78:@5157.4]
  assign _T_1888 = allocatedEntries_4 | initBits_4; // @[AxiLoadQueue.scala 73:78:@5158.4]
  assign _T_1889 = allocatedEntries_5 | initBits_5; // @[AxiLoadQueue.scala 73:78:@5159.4]
  assign _T_1890 = allocatedEntries_6 | initBits_6; // @[AxiLoadQueue.scala 73:78:@5160.4]
  assign _T_1891 = allocatedEntries_7 | initBits_7; // @[AxiLoadQueue.scala 73:78:@5161.4]
  assign _T_1892 = allocatedEntries_8 | initBits_8; // @[AxiLoadQueue.scala 73:78:@5162.4]
  assign _T_1893 = allocatedEntries_9 | initBits_9; // @[AxiLoadQueue.scala 73:78:@5163.4]
  assign _T_1894 = allocatedEntries_10 | initBits_10; // @[AxiLoadQueue.scala 73:78:@5164.4]
  assign _T_1895 = allocatedEntries_11 | initBits_11; // @[AxiLoadQueue.scala 73:78:@5165.4]
  assign _T_1896 = allocatedEntries_12 | initBits_12; // @[AxiLoadQueue.scala 73:78:@5166.4]
  assign _T_1897 = allocatedEntries_13 | initBits_13; // @[AxiLoadQueue.scala 73:78:@5167.4]
  assign _T_1898 = allocatedEntries_14 | initBits_14; // @[AxiLoadQueue.scala 73:78:@5168.4]
  assign _T_1899 = allocatedEntries_15 | initBits_15; // @[AxiLoadQueue.scala 73:78:@5169.4]
  assign _T_1930 = _T_1725[3:0]; // @[:@5209.6]
  assign _GEN_1 = 4'h1 == _T_1930 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_2 = 4'h2 == _T_1930 ? io_bbLoadOffsets_2 : _GEN_1; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_3 = 4'h3 == _T_1930 ? io_bbLoadOffsets_3 : _GEN_2; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_4 = 4'h4 == _T_1930 ? io_bbLoadOffsets_4 : _GEN_3; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_5 = 4'h5 == _T_1930 ? io_bbLoadOffsets_5 : _GEN_4; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_6 = 4'h6 == _T_1930 ? io_bbLoadOffsets_6 : _GEN_5; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_7 = 4'h7 == _T_1930 ? io_bbLoadOffsets_7 : _GEN_6; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_8 = 4'h8 == _T_1930 ? io_bbLoadOffsets_8 : _GEN_7; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_9 = 4'h9 == _T_1930 ? io_bbLoadOffsets_9 : _GEN_8; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_10 = 4'ha == _T_1930 ? io_bbLoadOffsets_10 : _GEN_9; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_11 = 4'hb == _T_1930 ? io_bbLoadOffsets_11 : _GEN_10; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_12 = 4'hc == _T_1930 ? io_bbLoadOffsets_12 : _GEN_11; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_13 = 4'hd == _T_1930 ? io_bbLoadOffsets_13 : _GEN_12; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_14 = 4'he == _T_1930 ? io_bbLoadOffsets_14 : _GEN_13; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_15 = 4'hf == _T_1930 ? io_bbLoadOffsets_15 : _GEN_14; // @[AxiLoadQueue.scala 77:20:@5210.6]
  assign _GEN_32 = initBits_0 ? _GEN_15 : offsetQ_0; // @[AxiLoadQueue.scala 76:25:@5203.4]
  assign _GEN_33 = initBits_0 ? 1'h0 : portQ_0; // @[AxiLoadQueue.scala 76:25:@5203.4]
  assign _T_1948 = _T_1734[3:0]; // @[:@5225.6]
  assign _GEN_35 = 4'h1 == _T_1948 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_36 = 4'h2 == _T_1948 ? io_bbLoadOffsets_2 : _GEN_35; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_37 = 4'h3 == _T_1948 ? io_bbLoadOffsets_3 : _GEN_36; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_38 = 4'h4 == _T_1948 ? io_bbLoadOffsets_4 : _GEN_37; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_39 = 4'h5 == _T_1948 ? io_bbLoadOffsets_5 : _GEN_38; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_40 = 4'h6 == _T_1948 ? io_bbLoadOffsets_6 : _GEN_39; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_41 = 4'h7 == _T_1948 ? io_bbLoadOffsets_7 : _GEN_40; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_42 = 4'h8 == _T_1948 ? io_bbLoadOffsets_8 : _GEN_41; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_43 = 4'h9 == _T_1948 ? io_bbLoadOffsets_9 : _GEN_42; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_44 = 4'ha == _T_1948 ? io_bbLoadOffsets_10 : _GEN_43; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_45 = 4'hb == _T_1948 ? io_bbLoadOffsets_11 : _GEN_44; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_46 = 4'hc == _T_1948 ? io_bbLoadOffsets_12 : _GEN_45; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_47 = 4'hd == _T_1948 ? io_bbLoadOffsets_13 : _GEN_46; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_48 = 4'he == _T_1948 ? io_bbLoadOffsets_14 : _GEN_47; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_49 = 4'hf == _T_1948 ? io_bbLoadOffsets_15 : _GEN_48; // @[AxiLoadQueue.scala 77:20:@5226.6]
  assign _GEN_66 = initBits_1 ? _GEN_49 : offsetQ_1; // @[AxiLoadQueue.scala 76:25:@5219.4]
  assign _GEN_67 = initBits_1 ? 1'h0 : portQ_1; // @[AxiLoadQueue.scala 76:25:@5219.4]
  assign _T_1966 = _T_1743[3:0]; // @[:@5241.6]
  assign _GEN_69 = 4'h1 == _T_1966 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_70 = 4'h2 == _T_1966 ? io_bbLoadOffsets_2 : _GEN_69; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_71 = 4'h3 == _T_1966 ? io_bbLoadOffsets_3 : _GEN_70; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_72 = 4'h4 == _T_1966 ? io_bbLoadOffsets_4 : _GEN_71; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_73 = 4'h5 == _T_1966 ? io_bbLoadOffsets_5 : _GEN_72; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_74 = 4'h6 == _T_1966 ? io_bbLoadOffsets_6 : _GEN_73; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_75 = 4'h7 == _T_1966 ? io_bbLoadOffsets_7 : _GEN_74; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_76 = 4'h8 == _T_1966 ? io_bbLoadOffsets_8 : _GEN_75; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_77 = 4'h9 == _T_1966 ? io_bbLoadOffsets_9 : _GEN_76; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_78 = 4'ha == _T_1966 ? io_bbLoadOffsets_10 : _GEN_77; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_79 = 4'hb == _T_1966 ? io_bbLoadOffsets_11 : _GEN_78; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_80 = 4'hc == _T_1966 ? io_bbLoadOffsets_12 : _GEN_79; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_81 = 4'hd == _T_1966 ? io_bbLoadOffsets_13 : _GEN_80; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_82 = 4'he == _T_1966 ? io_bbLoadOffsets_14 : _GEN_81; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_83 = 4'hf == _T_1966 ? io_bbLoadOffsets_15 : _GEN_82; // @[AxiLoadQueue.scala 77:20:@5242.6]
  assign _GEN_100 = initBits_2 ? _GEN_83 : offsetQ_2; // @[AxiLoadQueue.scala 76:25:@5235.4]
  assign _GEN_101 = initBits_2 ? 1'h0 : portQ_2; // @[AxiLoadQueue.scala 76:25:@5235.4]
  assign _T_1984 = _T_1752[3:0]; // @[:@5257.6]
  assign _GEN_103 = 4'h1 == _T_1984 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_104 = 4'h2 == _T_1984 ? io_bbLoadOffsets_2 : _GEN_103; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_105 = 4'h3 == _T_1984 ? io_bbLoadOffsets_3 : _GEN_104; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_106 = 4'h4 == _T_1984 ? io_bbLoadOffsets_4 : _GEN_105; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_107 = 4'h5 == _T_1984 ? io_bbLoadOffsets_5 : _GEN_106; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_108 = 4'h6 == _T_1984 ? io_bbLoadOffsets_6 : _GEN_107; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_109 = 4'h7 == _T_1984 ? io_bbLoadOffsets_7 : _GEN_108; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_110 = 4'h8 == _T_1984 ? io_bbLoadOffsets_8 : _GEN_109; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_111 = 4'h9 == _T_1984 ? io_bbLoadOffsets_9 : _GEN_110; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_112 = 4'ha == _T_1984 ? io_bbLoadOffsets_10 : _GEN_111; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_113 = 4'hb == _T_1984 ? io_bbLoadOffsets_11 : _GEN_112; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_114 = 4'hc == _T_1984 ? io_bbLoadOffsets_12 : _GEN_113; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_115 = 4'hd == _T_1984 ? io_bbLoadOffsets_13 : _GEN_114; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_116 = 4'he == _T_1984 ? io_bbLoadOffsets_14 : _GEN_115; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_117 = 4'hf == _T_1984 ? io_bbLoadOffsets_15 : _GEN_116; // @[AxiLoadQueue.scala 77:20:@5258.6]
  assign _GEN_134 = initBits_3 ? _GEN_117 : offsetQ_3; // @[AxiLoadQueue.scala 76:25:@5251.4]
  assign _GEN_135 = initBits_3 ? 1'h0 : portQ_3; // @[AxiLoadQueue.scala 76:25:@5251.4]
  assign _T_2002 = _T_1761[3:0]; // @[:@5273.6]
  assign _GEN_137 = 4'h1 == _T_2002 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_138 = 4'h2 == _T_2002 ? io_bbLoadOffsets_2 : _GEN_137; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_139 = 4'h3 == _T_2002 ? io_bbLoadOffsets_3 : _GEN_138; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_140 = 4'h4 == _T_2002 ? io_bbLoadOffsets_4 : _GEN_139; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_141 = 4'h5 == _T_2002 ? io_bbLoadOffsets_5 : _GEN_140; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_142 = 4'h6 == _T_2002 ? io_bbLoadOffsets_6 : _GEN_141; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_143 = 4'h7 == _T_2002 ? io_bbLoadOffsets_7 : _GEN_142; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_144 = 4'h8 == _T_2002 ? io_bbLoadOffsets_8 : _GEN_143; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_145 = 4'h9 == _T_2002 ? io_bbLoadOffsets_9 : _GEN_144; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_146 = 4'ha == _T_2002 ? io_bbLoadOffsets_10 : _GEN_145; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_147 = 4'hb == _T_2002 ? io_bbLoadOffsets_11 : _GEN_146; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_148 = 4'hc == _T_2002 ? io_bbLoadOffsets_12 : _GEN_147; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_149 = 4'hd == _T_2002 ? io_bbLoadOffsets_13 : _GEN_148; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_150 = 4'he == _T_2002 ? io_bbLoadOffsets_14 : _GEN_149; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_151 = 4'hf == _T_2002 ? io_bbLoadOffsets_15 : _GEN_150; // @[AxiLoadQueue.scala 77:20:@5274.6]
  assign _GEN_168 = initBits_4 ? _GEN_151 : offsetQ_4; // @[AxiLoadQueue.scala 76:25:@5267.4]
  assign _GEN_169 = initBits_4 ? 1'h0 : portQ_4; // @[AxiLoadQueue.scala 76:25:@5267.4]
  assign _T_2020 = _T_1770[3:0]; // @[:@5289.6]
  assign _GEN_171 = 4'h1 == _T_2020 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_172 = 4'h2 == _T_2020 ? io_bbLoadOffsets_2 : _GEN_171; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_173 = 4'h3 == _T_2020 ? io_bbLoadOffsets_3 : _GEN_172; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_174 = 4'h4 == _T_2020 ? io_bbLoadOffsets_4 : _GEN_173; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_175 = 4'h5 == _T_2020 ? io_bbLoadOffsets_5 : _GEN_174; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_176 = 4'h6 == _T_2020 ? io_bbLoadOffsets_6 : _GEN_175; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_177 = 4'h7 == _T_2020 ? io_bbLoadOffsets_7 : _GEN_176; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_178 = 4'h8 == _T_2020 ? io_bbLoadOffsets_8 : _GEN_177; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_179 = 4'h9 == _T_2020 ? io_bbLoadOffsets_9 : _GEN_178; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_180 = 4'ha == _T_2020 ? io_bbLoadOffsets_10 : _GEN_179; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_181 = 4'hb == _T_2020 ? io_bbLoadOffsets_11 : _GEN_180; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_182 = 4'hc == _T_2020 ? io_bbLoadOffsets_12 : _GEN_181; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_183 = 4'hd == _T_2020 ? io_bbLoadOffsets_13 : _GEN_182; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_184 = 4'he == _T_2020 ? io_bbLoadOffsets_14 : _GEN_183; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_185 = 4'hf == _T_2020 ? io_bbLoadOffsets_15 : _GEN_184; // @[AxiLoadQueue.scala 77:20:@5290.6]
  assign _GEN_202 = initBits_5 ? _GEN_185 : offsetQ_5; // @[AxiLoadQueue.scala 76:25:@5283.4]
  assign _GEN_203 = initBits_5 ? 1'h0 : portQ_5; // @[AxiLoadQueue.scala 76:25:@5283.4]
  assign _T_2038 = _T_1779[3:0]; // @[:@5305.6]
  assign _GEN_205 = 4'h1 == _T_2038 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_206 = 4'h2 == _T_2038 ? io_bbLoadOffsets_2 : _GEN_205; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_207 = 4'h3 == _T_2038 ? io_bbLoadOffsets_3 : _GEN_206; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_208 = 4'h4 == _T_2038 ? io_bbLoadOffsets_4 : _GEN_207; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_209 = 4'h5 == _T_2038 ? io_bbLoadOffsets_5 : _GEN_208; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_210 = 4'h6 == _T_2038 ? io_bbLoadOffsets_6 : _GEN_209; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_211 = 4'h7 == _T_2038 ? io_bbLoadOffsets_7 : _GEN_210; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_212 = 4'h8 == _T_2038 ? io_bbLoadOffsets_8 : _GEN_211; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_213 = 4'h9 == _T_2038 ? io_bbLoadOffsets_9 : _GEN_212; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_214 = 4'ha == _T_2038 ? io_bbLoadOffsets_10 : _GEN_213; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_215 = 4'hb == _T_2038 ? io_bbLoadOffsets_11 : _GEN_214; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_216 = 4'hc == _T_2038 ? io_bbLoadOffsets_12 : _GEN_215; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_217 = 4'hd == _T_2038 ? io_bbLoadOffsets_13 : _GEN_216; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_218 = 4'he == _T_2038 ? io_bbLoadOffsets_14 : _GEN_217; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_219 = 4'hf == _T_2038 ? io_bbLoadOffsets_15 : _GEN_218; // @[AxiLoadQueue.scala 77:20:@5306.6]
  assign _GEN_236 = initBits_6 ? _GEN_219 : offsetQ_6; // @[AxiLoadQueue.scala 76:25:@5299.4]
  assign _GEN_237 = initBits_6 ? 1'h0 : portQ_6; // @[AxiLoadQueue.scala 76:25:@5299.4]
  assign _T_2056 = _T_1788[3:0]; // @[:@5321.6]
  assign _GEN_239 = 4'h1 == _T_2056 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_240 = 4'h2 == _T_2056 ? io_bbLoadOffsets_2 : _GEN_239; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_241 = 4'h3 == _T_2056 ? io_bbLoadOffsets_3 : _GEN_240; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_242 = 4'h4 == _T_2056 ? io_bbLoadOffsets_4 : _GEN_241; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_243 = 4'h5 == _T_2056 ? io_bbLoadOffsets_5 : _GEN_242; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_244 = 4'h6 == _T_2056 ? io_bbLoadOffsets_6 : _GEN_243; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_245 = 4'h7 == _T_2056 ? io_bbLoadOffsets_7 : _GEN_244; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_246 = 4'h8 == _T_2056 ? io_bbLoadOffsets_8 : _GEN_245; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_247 = 4'h9 == _T_2056 ? io_bbLoadOffsets_9 : _GEN_246; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_248 = 4'ha == _T_2056 ? io_bbLoadOffsets_10 : _GEN_247; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_249 = 4'hb == _T_2056 ? io_bbLoadOffsets_11 : _GEN_248; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_250 = 4'hc == _T_2056 ? io_bbLoadOffsets_12 : _GEN_249; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_251 = 4'hd == _T_2056 ? io_bbLoadOffsets_13 : _GEN_250; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_252 = 4'he == _T_2056 ? io_bbLoadOffsets_14 : _GEN_251; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_253 = 4'hf == _T_2056 ? io_bbLoadOffsets_15 : _GEN_252; // @[AxiLoadQueue.scala 77:20:@5322.6]
  assign _GEN_270 = initBits_7 ? _GEN_253 : offsetQ_7; // @[AxiLoadQueue.scala 76:25:@5315.4]
  assign _GEN_271 = initBits_7 ? 1'h0 : portQ_7; // @[AxiLoadQueue.scala 76:25:@5315.4]
  assign _T_2074 = _T_1797[3:0]; // @[:@5337.6]
  assign _GEN_273 = 4'h1 == _T_2074 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_274 = 4'h2 == _T_2074 ? io_bbLoadOffsets_2 : _GEN_273; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_275 = 4'h3 == _T_2074 ? io_bbLoadOffsets_3 : _GEN_274; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_276 = 4'h4 == _T_2074 ? io_bbLoadOffsets_4 : _GEN_275; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_277 = 4'h5 == _T_2074 ? io_bbLoadOffsets_5 : _GEN_276; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_278 = 4'h6 == _T_2074 ? io_bbLoadOffsets_6 : _GEN_277; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_279 = 4'h7 == _T_2074 ? io_bbLoadOffsets_7 : _GEN_278; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_280 = 4'h8 == _T_2074 ? io_bbLoadOffsets_8 : _GEN_279; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_281 = 4'h9 == _T_2074 ? io_bbLoadOffsets_9 : _GEN_280; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_282 = 4'ha == _T_2074 ? io_bbLoadOffsets_10 : _GEN_281; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_283 = 4'hb == _T_2074 ? io_bbLoadOffsets_11 : _GEN_282; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_284 = 4'hc == _T_2074 ? io_bbLoadOffsets_12 : _GEN_283; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_285 = 4'hd == _T_2074 ? io_bbLoadOffsets_13 : _GEN_284; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_286 = 4'he == _T_2074 ? io_bbLoadOffsets_14 : _GEN_285; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_287 = 4'hf == _T_2074 ? io_bbLoadOffsets_15 : _GEN_286; // @[AxiLoadQueue.scala 77:20:@5338.6]
  assign _GEN_304 = initBits_8 ? _GEN_287 : offsetQ_8; // @[AxiLoadQueue.scala 76:25:@5331.4]
  assign _GEN_305 = initBits_8 ? 1'h0 : portQ_8; // @[AxiLoadQueue.scala 76:25:@5331.4]
  assign _T_2092 = _T_1806[3:0]; // @[:@5353.6]
  assign _GEN_307 = 4'h1 == _T_2092 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_308 = 4'h2 == _T_2092 ? io_bbLoadOffsets_2 : _GEN_307; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_309 = 4'h3 == _T_2092 ? io_bbLoadOffsets_3 : _GEN_308; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_310 = 4'h4 == _T_2092 ? io_bbLoadOffsets_4 : _GEN_309; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_311 = 4'h5 == _T_2092 ? io_bbLoadOffsets_5 : _GEN_310; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_312 = 4'h6 == _T_2092 ? io_bbLoadOffsets_6 : _GEN_311; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_313 = 4'h7 == _T_2092 ? io_bbLoadOffsets_7 : _GEN_312; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_314 = 4'h8 == _T_2092 ? io_bbLoadOffsets_8 : _GEN_313; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_315 = 4'h9 == _T_2092 ? io_bbLoadOffsets_9 : _GEN_314; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_316 = 4'ha == _T_2092 ? io_bbLoadOffsets_10 : _GEN_315; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_317 = 4'hb == _T_2092 ? io_bbLoadOffsets_11 : _GEN_316; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_318 = 4'hc == _T_2092 ? io_bbLoadOffsets_12 : _GEN_317; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_319 = 4'hd == _T_2092 ? io_bbLoadOffsets_13 : _GEN_318; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_320 = 4'he == _T_2092 ? io_bbLoadOffsets_14 : _GEN_319; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_321 = 4'hf == _T_2092 ? io_bbLoadOffsets_15 : _GEN_320; // @[AxiLoadQueue.scala 77:20:@5354.6]
  assign _GEN_338 = initBits_9 ? _GEN_321 : offsetQ_9; // @[AxiLoadQueue.scala 76:25:@5347.4]
  assign _GEN_339 = initBits_9 ? 1'h0 : portQ_9; // @[AxiLoadQueue.scala 76:25:@5347.4]
  assign _T_2110 = _T_1815[3:0]; // @[:@5369.6]
  assign _GEN_341 = 4'h1 == _T_2110 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_342 = 4'h2 == _T_2110 ? io_bbLoadOffsets_2 : _GEN_341; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_343 = 4'h3 == _T_2110 ? io_bbLoadOffsets_3 : _GEN_342; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_344 = 4'h4 == _T_2110 ? io_bbLoadOffsets_4 : _GEN_343; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_345 = 4'h5 == _T_2110 ? io_bbLoadOffsets_5 : _GEN_344; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_346 = 4'h6 == _T_2110 ? io_bbLoadOffsets_6 : _GEN_345; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_347 = 4'h7 == _T_2110 ? io_bbLoadOffsets_7 : _GEN_346; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_348 = 4'h8 == _T_2110 ? io_bbLoadOffsets_8 : _GEN_347; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_349 = 4'h9 == _T_2110 ? io_bbLoadOffsets_9 : _GEN_348; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_350 = 4'ha == _T_2110 ? io_bbLoadOffsets_10 : _GEN_349; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_351 = 4'hb == _T_2110 ? io_bbLoadOffsets_11 : _GEN_350; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_352 = 4'hc == _T_2110 ? io_bbLoadOffsets_12 : _GEN_351; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_353 = 4'hd == _T_2110 ? io_bbLoadOffsets_13 : _GEN_352; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_354 = 4'he == _T_2110 ? io_bbLoadOffsets_14 : _GEN_353; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_355 = 4'hf == _T_2110 ? io_bbLoadOffsets_15 : _GEN_354; // @[AxiLoadQueue.scala 77:20:@5370.6]
  assign _GEN_372 = initBits_10 ? _GEN_355 : offsetQ_10; // @[AxiLoadQueue.scala 76:25:@5363.4]
  assign _GEN_373 = initBits_10 ? 1'h0 : portQ_10; // @[AxiLoadQueue.scala 76:25:@5363.4]
  assign _T_2128 = _T_1824[3:0]; // @[:@5385.6]
  assign _GEN_375 = 4'h1 == _T_2128 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_376 = 4'h2 == _T_2128 ? io_bbLoadOffsets_2 : _GEN_375; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_377 = 4'h3 == _T_2128 ? io_bbLoadOffsets_3 : _GEN_376; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_378 = 4'h4 == _T_2128 ? io_bbLoadOffsets_4 : _GEN_377; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_379 = 4'h5 == _T_2128 ? io_bbLoadOffsets_5 : _GEN_378; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_380 = 4'h6 == _T_2128 ? io_bbLoadOffsets_6 : _GEN_379; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_381 = 4'h7 == _T_2128 ? io_bbLoadOffsets_7 : _GEN_380; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_382 = 4'h8 == _T_2128 ? io_bbLoadOffsets_8 : _GEN_381; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_383 = 4'h9 == _T_2128 ? io_bbLoadOffsets_9 : _GEN_382; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_384 = 4'ha == _T_2128 ? io_bbLoadOffsets_10 : _GEN_383; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_385 = 4'hb == _T_2128 ? io_bbLoadOffsets_11 : _GEN_384; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_386 = 4'hc == _T_2128 ? io_bbLoadOffsets_12 : _GEN_385; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_387 = 4'hd == _T_2128 ? io_bbLoadOffsets_13 : _GEN_386; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_388 = 4'he == _T_2128 ? io_bbLoadOffsets_14 : _GEN_387; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_389 = 4'hf == _T_2128 ? io_bbLoadOffsets_15 : _GEN_388; // @[AxiLoadQueue.scala 77:20:@5386.6]
  assign _GEN_406 = initBits_11 ? _GEN_389 : offsetQ_11; // @[AxiLoadQueue.scala 76:25:@5379.4]
  assign _GEN_407 = initBits_11 ? 1'h0 : portQ_11; // @[AxiLoadQueue.scala 76:25:@5379.4]
  assign _T_2146 = _T_1833[3:0]; // @[:@5401.6]
  assign _GEN_409 = 4'h1 == _T_2146 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_410 = 4'h2 == _T_2146 ? io_bbLoadOffsets_2 : _GEN_409; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_411 = 4'h3 == _T_2146 ? io_bbLoadOffsets_3 : _GEN_410; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_412 = 4'h4 == _T_2146 ? io_bbLoadOffsets_4 : _GEN_411; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_413 = 4'h5 == _T_2146 ? io_bbLoadOffsets_5 : _GEN_412; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_414 = 4'h6 == _T_2146 ? io_bbLoadOffsets_6 : _GEN_413; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_415 = 4'h7 == _T_2146 ? io_bbLoadOffsets_7 : _GEN_414; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_416 = 4'h8 == _T_2146 ? io_bbLoadOffsets_8 : _GEN_415; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_417 = 4'h9 == _T_2146 ? io_bbLoadOffsets_9 : _GEN_416; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_418 = 4'ha == _T_2146 ? io_bbLoadOffsets_10 : _GEN_417; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_419 = 4'hb == _T_2146 ? io_bbLoadOffsets_11 : _GEN_418; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_420 = 4'hc == _T_2146 ? io_bbLoadOffsets_12 : _GEN_419; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_421 = 4'hd == _T_2146 ? io_bbLoadOffsets_13 : _GEN_420; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_422 = 4'he == _T_2146 ? io_bbLoadOffsets_14 : _GEN_421; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_423 = 4'hf == _T_2146 ? io_bbLoadOffsets_15 : _GEN_422; // @[AxiLoadQueue.scala 77:20:@5402.6]
  assign _GEN_440 = initBits_12 ? _GEN_423 : offsetQ_12; // @[AxiLoadQueue.scala 76:25:@5395.4]
  assign _GEN_441 = initBits_12 ? 1'h0 : portQ_12; // @[AxiLoadQueue.scala 76:25:@5395.4]
  assign _T_2164 = _T_1842[3:0]; // @[:@5417.6]
  assign _GEN_443 = 4'h1 == _T_2164 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_444 = 4'h2 == _T_2164 ? io_bbLoadOffsets_2 : _GEN_443; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_445 = 4'h3 == _T_2164 ? io_bbLoadOffsets_3 : _GEN_444; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_446 = 4'h4 == _T_2164 ? io_bbLoadOffsets_4 : _GEN_445; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_447 = 4'h5 == _T_2164 ? io_bbLoadOffsets_5 : _GEN_446; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_448 = 4'h6 == _T_2164 ? io_bbLoadOffsets_6 : _GEN_447; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_449 = 4'h7 == _T_2164 ? io_bbLoadOffsets_7 : _GEN_448; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_450 = 4'h8 == _T_2164 ? io_bbLoadOffsets_8 : _GEN_449; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_451 = 4'h9 == _T_2164 ? io_bbLoadOffsets_9 : _GEN_450; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_452 = 4'ha == _T_2164 ? io_bbLoadOffsets_10 : _GEN_451; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_453 = 4'hb == _T_2164 ? io_bbLoadOffsets_11 : _GEN_452; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_454 = 4'hc == _T_2164 ? io_bbLoadOffsets_12 : _GEN_453; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_455 = 4'hd == _T_2164 ? io_bbLoadOffsets_13 : _GEN_454; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_456 = 4'he == _T_2164 ? io_bbLoadOffsets_14 : _GEN_455; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_457 = 4'hf == _T_2164 ? io_bbLoadOffsets_15 : _GEN_456; // @[AxiLoadQueue.scala 77:20:@5418.6]
  assign _GEN_474 = initBits_13 ? _GEN_457 : offsetQ_13; // @[AxiLoadQueue.scala 76:25:@5411.4]
  assign _GEN_475 = initBits_13 ? 1'h0 : portQ_13; // @[AxiLoadQueue.scala 76:25:@5411.4]
  assign _T_2182 = _T_1851[3:0]; // @[:@5433.6]
  assign _GEN_477 = 4'h1 == _T_2182 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_478 = 4'h2 == _T_2182 ? io_bbLoadOffsets_2 : _GEN_477; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_479 = 4'h3 == _T_2182 ? io_bbLoadOffsets_3 : _GEN_478; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_480 = 4'h4 == _T_2182 ? io_bbLoadOffsets_4 : _GEN_479; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_481 = 4'h5 == _T_2182 ? io_bbLoadOffsets_5 : _GEN_480; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_482 = 4'h6 == _T_2182 ? io_bbLoadOffsets_6 : _GEN_481; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_483 = 4'h7 == _T_2182 ? io_bbLoadOffsets_7 : _GEN_482; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_484 = 4'h8 == _T_2182 ? io_bbLoadOffsets_8 : _GEN_483; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_485 = 4'h9 == _T_2182 ? io_bbLoadOffsets_9 : _GEN_484; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_486 = 4'ha == _T_2182 ? io_bbLoadOffsets_10 : _GEN_485; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_487 = 4'hb == _T_2182 ? io_bbLoadOffsets_11 : _GEN_486; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_488 = 4'hc == _T_2182 ? io_bbLoadOffsets_12 : _GEN_487; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_489 = 4'hd == _T_2182 ? io_bbLoadOffsets_13 : _GEN_488; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_490 = 4'he == _T_2182 ? io_bbLoadOffsets_14 : _GEN_489; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_491 = 4'hf == _T_2182 ? io_bbLoadOffsets_15 : _GEN_490; // @[AxiLoadQueue.scala 77:20:@5434.6]
  assign _GEN_508 = initBits_14 ? _GEN_491 : offsetQ_14; // @[AxiLoadQueue.scala 76:25:@5427.4]
  assign _GEN_509 = initBits_14 ? 1'h0 : portQ_14; // @[AxiLoadQueue.scala 76:25:@5427.4]
  assign _T_2200 = _T_1860[3:0]; // @[:@5449.6]
  assign _GEN_511 = 4'h1 == _T_2200 ? io_bbLoadOffsets_1 : io_bbLoadOffsets_0; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_512 = 4'h2 == _T_2200 ? io_bbLoadOffsets_2 : _GEN_511; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_513 = 4'h3 == _T_2200 ? io_bbLoadOffsets_3 : _GEN_512; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_514 = 4'h4 == _T_2200 ? io_bbLoadOffsets_4 : _GEN_513; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_515 = 4'h5 == _T_2200 ? io_bbLoadOffsets_5 : _GEN_514; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_516 = 4'h6 == _T_2200 ? io_bbLoadOffsets_6 : _GEN_515; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_517 = 4'h7 == _T_2200 ? io_bbLoadOffsets_7 : _GEN_516; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_518 = 4'h8 == _T_2200 ? io_bbLoadOffsets_8 : _GEN_517; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_519 = 4'h9 == _T_2200 ? io_bbLoadOffsets_9 : _GEN_518; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_520 = 4'ha == _T_2200 ? io_bbLoadOffsets_10 : _GEN_519; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_521 = 4'hb == _T_2200 ? io_bbLoadOffsets_11 : _GEN_520; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_522 = 4'hc == _T_2200 ? io_bbLoadOffsets_12 : _GEN_521; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_523 = 4'hd == _T_2200 ? io_bbLoadOffsets_13 : _GEN_522; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_524 = 4'he == _T_2200 ? io_bbLoadOffsets_14 : _GEN_523; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_525 = 4'hf == _T_2200 ? io_bbLoadOffsets_15 : _GEN_524; // @[AxiLoadQueue.scala 77:20:@5450.6]
  assign _GEN_542 = initBits_15 ? _GEN_525 : offsetQ_15; // @[AxiLoadQueue.scala 76:25:@5443.4]
  assign _GEN_543 = initBits_15 ? 1'h0 : portQ_15; // @[AxiLoadQueue.scala 76:25:@5443.4]
  assign _T_2222 = _GEN_15 + 4'h1; // @[util.scala 10:8:@5468.6]
  assign _GEN_31 = _T_2222 % 5'h10; // @[util.scala 10:14:@5469.6]
  assign _T_2223 = _GEN_31[4:0]; // @[util.scala 10:14:@5469.6]
  assign _GEN_2341 = {{1'd0}, io_storeTail}; // @[AxiLoadQueue.scala 97:56:@5470.6]
  assign _T_2224 = _T_2223 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5470.6]
  assign _T_2225 = io_storeEmpty & _T_2224; // @[AxiLoadQueue.scala 96:50:@5471.6]
  assign _T_2227 = _T_2225 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5472.6]
  assign _T_2229 = previousStoreHead <= offsetQ_0; // @[AxiLoadQueue.scala 101:36:@5480.8]
  assign _T_2230 = offsetQ_0 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5481.8]
  assign _T_2231 = _T_2229 & _T_2230; // @[AxiLoadQueue.scala 101:61:@5482.8]
  assign _T_2233 = previousStoreHead > io_storeHead; // @[AxiLoadQueue.scala 103:36:@5487.10]
  assign _T_2234 = io_storeHead <= offsetQ_0; // @[AxiLoadQueue.scala 103:69:@5488.10]
  assign _T_2235 = offsetQ_0 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5489.10]
  assign _T_2236 = _T_2234 & _T_2235; // @[AxiLoadQueue.scala 103:94:@5490.10]
  assign _T_2238 = _T_2236 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5491.10]
  assign _T_2239 = _T_2233 & _T_2238; // @[AxiLoadQueue.scala 103:51:@5492.10]
  assign _GEN_560 = _T_2239 ? 1'h0 : checkBits_0; // @[AxiLoadQueue.scala 104:53:@5493.10]
  assign _GEN_561 = _T_2231 ? 1'h0 : _GEN_560; // @[AxiLoadQueue.scala 101:102:@5483.8]
  assign _GEN_562 = io_storeEmpty ? 1'h0 : _GEN_561; // @[AxiLoadQueue.scala 99:27:@5476.6]
  assign _GEN_563 = initBits_0 ? _T_2227 : _GEN_562; // @[AxiLoadQueue.scala 95:34:@5461.4]
  assign _T_2252 = _GEN_49 + 4'h1; // @[util.scala 10:8:@5504.6]
  assign _GEN_34 = _T_2252 % 5'h10; // @[util.scala 10:14:@5505.6]
  assign _T_2253 = _GEN_34[4:0]; // @[util.scala 10:14:@5505.6]
  assign _T_2254 = _T_2253 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5506.6]
  assign _T_2255 = io_storeEmpty & _T_2254; // @[AxiLoadQueue.scala 96:50:@5507.6]
  assign _T_2257 = _T_2255 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5508.6]
  assign _T_2259 = previousStoreHead <= offsetQ_1; // @[AxiLoadQueue.scala 101:36:@5516.8]
  assign _T_2260 = offsetQ_1 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5517.8]
  assign _T_2261 = _T_2259 & _T_2260; // @[AxiLoadQueue.scala 101:61:@5518.8]
  assign _T_2264 = io_storeHead <= offsetQ_1; // @[AxiLoadQueue.scala 103:69:@5524.10]
  assign _T_2265 = offsetQ_1 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5525.10]
  assign _T_2266 = _T_2264 & _T_2265; // @[AxiLoadQueue.scala 103:94:@5526.10]
  assign _T_2268 = _T_2266 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5527.10]
  assign _T_2269 = _T_2233 & _T_2268; // @[AxiLoadQueue.scala 103:51:@5528.10]
  assign _GEN_580 = _T_2269 ? 1'h0 : checkBits_1; // @[AxiLoadQueue.scala 104:53:@5529.10]
  assign _GEN_581 = _T_2261 ? 1'h0 : _GEN_580; // @[AxiLoadQueue.scala 101:102:@5519.8]
  assign _GEN_582 = io_storeEmpty ? 1'h0 : _GEN_581; // @[AxiLoadQueue.scala 99:27:@5512.6]
  assign _GEN_583 = initBits_1 ? _T_2257 : _GEN_582; // @[AxiLoadQueue.scala 95:34:@5497.4]
  assign _T_2282 = _GEN_83 + 4'h1; // @[util.scala 10:8:@5540.6]
  assign _GEN_50 = _T_2282 % 5'h10; // @[util.scala 10:14:@5541.6]
  assign _T_2283 = _GEN_50[4:0]; // @[util.scala 10:14:@5541.6]
  assign _T_2284 = _T_2283 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5542.6]
  assign _T_2285 = io_storeEmpty & _T_2284; // @[AxiLoadQueue.scala 96:50:@5543.6]
  assign _T_2287 = _T_2285 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5544.6]
  assign _T_2289 = previousStoreHead <= offsetQ_2; // @[AxiLoadQueue.scala 101:36:@5552.8]
  assign _T_2290 = offsetQ_2 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5553.8]
  assign _T_2291 = _T_2289 & _T_2290; // @[AxiLoadQueue.scala 101:61:@5554.8]
  assign _T_2294 = io_storeHead <= offsetQ_2; // @[AxiLoadQueue.scala 103:69:@5560.10]
  assign _T_2295 = offsetQ_2 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5561.10]
  assign _T_2296 = _T_2294 & _T_2295; // @[AxiLoadQueue.scala 103:94:@5562.10]
  assign _T_2298 = _T_2296 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5563.10]
  assign _T_2299 = _T_2233 & _T_2298; // @[AxiLoadQueue.scala 103:51:@5564.10]
  assign _GEN_600 = _T_2299 ? 1'h0 : checkBits_2; // @[AxiLoadQueue.scala 104:53:@5565.10]
  assign _GEN_601 = _T_2291 ? 1'h0 : _GEN_600; // @[AxiLoadQueue.scala 101:102:@5555.8]
  assign _GEN_602 = io_storeEmpty ? 1'h0 : _GEN_601; // @[AxiLoadQueue.scala 99:27:@5548.6]
  assign _GEN_603 = initBits_2 ? _T_2287 : _GEN_602; // @[AxiLoadQueue.scala 95:34:@5533.4]
  assign _T_2312 = _GEN_117 + 4'h1; // @[util.scala 10:8:@5576.6]
  assign _GEN_51 = _T_2312 % 5'h10; // @[util.scala 10:14:@5577.6]
  assign _T_2313 = _GEN_51[4:0]; // @[util.scala 10:14:@5577.6]
  assign _T_2314 = _T_2313 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5578.6]
  assign _T_2315 = io_storeEmpty & _T_2314; // @[AxiLoadQueue.scala 96:50:@5579.6]
  assign _T_2317 = _T_2315 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5580.6]
  assign _T_2319 = previousStoreHead <= offsetQ_3; // @[AxiLoadQueue.scala 101:36:@5588.8]
  assign _T_2320 = offsetQ_3 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5589.8]
  assign _T_2321 = _T_2319 & _T_2320; // @[AxiLoadQueue.scala 101:61:@5590.8]
  assign _T_2324 = io_storeHead <= offsetQ_3; // @[AxiLoadQueue.scala 103:69:@5596.10]
  assign _T_2325 = offsetQ_3 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5597.10]
  assign _T_2326 = _T_2324 & _T_2325; // @[AxiLoadQueue.scala 103:94:@5598.10]
  assign _T_2328 = _T_2326 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5599.10]
  assign _T_2329 = _T_2233 & _T_2328; // @[AxiLoadQueue.scala 103:51:@5600.10]
  assign _GEN_620 = _T_2329 ? 1'h0 : checkBits_3; // @[AxiLoadQueue.scala 104:53:@5601.10]
  assign _GEN_621 = _T_2321 ? 1'h0 : _GEN_620; // @[AxiLoadQueue.scala 101:102:@5591.8]
  assign _GEN_622 = io_storeEmpty ? 1'h0 : _GEN_621; // @[AxiLoadQueue.scala 99:27:@5584.6]
  assign _GEN_623 = initBits_3 ? _T_2317 : _GEN_622; // @[AxiLoadQueue.scala 95:34:@5569.4]
  assign _T_2342 = _GEN_151 + 4'h1; // @[util.scala 10:8:@5612.6]
  assign _GEN_52 = _T_2342 % 5'h10; // @[util.scala 10:14:@5613.6]
  assign _T_2343 = _GEN_52[4:0]; // @[util.scala 10:14:@5613.6]
  assign _T_2344 = _T_2343 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5614.6]
  assign _T_2345 = io_storeEmpty & _T_2344; // @[AxiLoadQueue.scala 96:50:@5615.6]
  assign _T_2347 = _T_2345 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5616.6]
  assign _T_2349 = previousStoreHead <= offsetQ_4; // @[AxiLoadQueue.scala 101:36:@5624.8]
  assign _T_2350 = offsetQ_4 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5625.8]
  assign _T_2351 = _T_2349 & _T_2350; // @[AxiLoadQueue.scala 101:61:@5626.8]
  assign _T_2354 = io_storeHead <= offsetQ_4; // @[AxiLoadQueue.scala 103:69:@5632.10]
  assign _T_2355 = offsetQ_4 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5633.10]
  assign _T_2356 = _T_2354 & _T_2355; // @[AxiLoadQueue.scala 103:94:@5634.10]
  assign _T_2358 = _T_2356 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5635.10]
  assign _T_2359 = _T_2233 & _T_2358; // @[AxiLoadQueue.scala 103:51:@5636.10]
  assign _GEN_640 = _T_2359 ? 1'h0 : checkBits_4; // @[AxiLoadQueue.scala 104:53:@5637.10]
  assign _GEN_641 = _T_2351 ? 1'h0 : _GEN_640; // @[AxiLoadQueue.scala 101:102:@5627.8]
  assign _GEN_642 = io_storeEmpty ? 1'h0 : _GEN_641; // @[AxiLoadQueue.scala 99:27:@5620.6]
  assign _GEN_643 = initBits_4 ? _T_2347 : _GEN_642; // @[AxiLoadQueue.scala 95:34:@5605.4]
  assign _T_2372 = _GEN_185 + 4'h1; // @[util.scala 10:8:@5648.6]
  assign _GEN_53 = _T_2372 % 5'h10; // @[util.scala 10:14:@5649.6]
  assign _T_2373 = _GEN_53[4:0]; // @[util.scala 10:14:@5649.6]
  assign _T_2374 = _T_2373 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5650.6]
  assign _T_2375 = io_storeEmpty & _T_2374; // @[AxiLoadQueue.scala 96:50:@5651.6]
  assign _T_2377 = _T_2375 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5652.6]
  assign _T_2379 = previousStoreHead <= offsetQ_5; // @[AxiLoadQueue.scala 101:36:@5660.8]
  assign _T_2380 = offsetQ_5 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5661.8]
  assign _T_2381 = _T_2379 & _T_2380; // @[AxiLoadQueue.scala 101:61:@5662.8]
  assign _T_2384 = io_storeHead <= offsetQ_5; // @[AxiLoadQueue.scala 103:69:@5668.10]
  assign _T_2385 = offsetQ_5 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5669.10]
  assign _T_2386 = _T_2384 & _T_2385; // @[AxiLoadQueue.scala 103:94:@5670.10]
  assign _T_2388 = _T_2386 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5671.10]
  assign _T_2389 = _T_2233 & _T_2388; // @[AxiLoadQueue.scala 103:51:@5672.10]
  assign _GEN_660 = _T_2389 ? 1'h0 : checkBits_5; // @[AxiLoadQueue.scala 104:53:@5673.10]
  assign _GEN_661 = _T_2381 ? 1'h0 : _GEN_660; // @[AxiLoadQueue.scala 101:102:@5663.8]
  assign _GEN_662 = io_storeEmpty ? 1'h0 : _GEN_661; // @[AxiLoadQueue.scala 99:27:@5656.6]
  assign _GEN_663 = initBits_5 ? _T_2377 : _GEN_662; // @[AxiLoadQueue.scala 95:34:@5641.4]
  assign _T_2402 = _GEN_219 + 4'h1; // @[util.scala 10:8:@5684.6]
  assign _GEN_54 = _T_2402 % 5'h10; // @[util.scala 10:14:@5685.6]
  assign _T_2403 = _GEN_54[4:0]; // @[util.scala 10:14:@5685.6]
  assign _T_2404 = _T_2403 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5686.6]
  assign _T_2405 = io_storeEmpty & _T_2404; // @[AxiLoadQueue.scala 96:50:@5687.6]
  assign _T_2407 = _T_2405 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5688.6]
  assign _T_2409 = previousStoreHead <= offsetQ_6; // @[AxiLoadQueue.scala 101:36:@5696.8]
  assign _T_2410 = offsetQ_6 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5697.8]
  assign _T_2411 = _T_2409 & _T_2410; // @[AxiLoadQueue.scala 101:61:@5698.8]
  assign _T_2414 = io_storeHead <= offsetQ_6; // @[AxiLoadQueue.scala 103:69:@5704.10]
  assign _T_2415 = offsetQ_6 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5705.10]
  assign _T_2416 = _T_2414 & _T_2415; // @[AxiLoadQueue.scala 103:94:@5706.10]
  assign _T_2418 = _T_2416 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5707.10]
  assign _T_2419 = _T_2233 & _T_2418; // @[AxiLoadQueue.scala 103:51:@5708.10]
  assign _GEN_680 = _T_2419 ? 1'h0 : checkBits_6; // @[AxiLoadQueue.scala 104:53:@5709.10]
  assign _GEN_681 = _T_2411 ? 1'h0 : _GEN_680; // @[AxiLoadQueue.scala 101:102:@5699.8]
  assign _GEN_682 = io_storeEmpty ? 1'h0 : _GEN_681; // @[AxiLoadQueue.scala 99:27:@5692.6]
  assign _GEN_683 = initBits_6 ? _T_2407 : _GEN_682; // @[AxiLoadQueue.scala 95:34:@5677.4]
  assign _T_2432 = _GEN_253 + 4'h1; // @[util.scala 10:8:@5720.6]
  assign _GEN_55 = _T_2432 % 5'h10; // @[util.scala 10:14:@5721.6]
  assign _T_2433 = _GEN_55[4:0]; // @[util.scala 10:14:@5721.6]
  assign _T_2434 = _T_2433 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5722.6]
  assign _T_2435 = io_storeEmpty & _T_2434; // @[AxiLoadQueue.scala 96:50:@5723.6]
  assign _T_2437 = _T_2435 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5724.6]
  assign _T_2439 = previousStoreHead <= offsetQ_7; // @[AxiLoadQueue.scala 101:36:@5732.8]
  assign _T_2440 = offsetQ_7 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5733.8]
  assign _T_2441 = _T_2439 & _T_2440; // @[AxiLoadQueue.scala 101:61:@5734.8]
  assign _T_2444 = io_storeHead <= offsetQ_7; // @[AxiLoadQueue.scala 103:69:@5740.10]
  assign _T_2445 = offsetQ_7 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5741.10]
  assign _T_2446 = _T_2444 & _T_2445; // @[AxiLoadQueue.scala 103:94:@5742.10]
  assign _T_2448 = _T_2446 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5743.10]
  assign _T_2449 = _T_2233 & _T_2448; // @[AxiLoadQueue.scala 103:51:@5744.10]
  assign _GEN_700 = _T_2449 ? 1'h0 : checkBits_7; // @[AxiLoadQueue.scala 104:53:@5745.10]
  assign _GEN_701 = _T_2441 ? 1'h0 : _GEN_700; // @[AxiLoadQueue.scala 101:102:@5735.8]
  assign _GEN_702 = io_storeEmpty ? 1'h0 : _GEN_701; // @[AxiLoadQueue.scala 99:27:@5728.6]
  assign _GEN_703 = initBits_7 ? _T_2437 : _GEN_702; // @[AxiLoadQueue.scala 95:34:@5713.4]
  assign _T_2462 = _GEN_287 + 4'h1; // @[util.scala 10:8:@5756.6]
  assign _GEN_56 = _T_2462 % 5'h10; // @[util.scala 10:14:@5757.6]
  assign _T_2463 = _GEN_56[4:0]; // @[util.scala 10:14:@5757.6]
  assign _T_2464 = _T_2463 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5758.6]
  assign _T_2465 = io_storeEmpty & _T_2464; // @[AxiLoadQueue.scala 96:50:@5759.6]
  assign _T_2467 = _T_2465 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5760.6]
  assign _T_2469 = previousStoreHead <= offsetQ_8; // @[AxiLoadQueue.scala 101:36:@5768.8]
  assign _T_2470 = offsetQ_8 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5769.8]
  assign _T_2471 = _T_2469 & _T_2470; // @[AxiLoadQueue.scala 101:61:@5770.8]
  assign _T_2474 = io_storeHead <= offsetQ_8; // @[AxiLoadQueue.scala 103:69:@5776.10]
  assign _T_2475 = offsetQ_8 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5777.10]
  assign _T_2476 = _T_2474 & _T_2475; // @[AxiLoadQueue.scala 103:94:@5778.10]
  assign _T_2478 = _T_2476 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5779.10]
  assign _T_2479 = _T_2233 & _T_2478; // @[AxiLoadQueue.scala 103:51:@5780.10]
  assign _GEN_720 = _T_2479 ? 1'h0 : checkBits_8; // @[AxiLoadQueue.scala 104:53:@5781.10]
  assign _GEN_721 = _T_2471 ? 1'h0 : _GEN_720; // @[AxiLoadQueue.scala 101:102:@5771.8]
  assign _GEN_722 = io_storeEmpty ? 1'h0 : _GEN_721; // @[AxiLoadQueue.scala 99:27:@5764.6]
  assign _GEN_723 = initBits_8 ? _T_2467 : _GEN_722; // @[AxiLoadQueue.scala 95:34:@5749.4]
  assign _T_2492 = _GEN_321 + 4'h1; // @[util.scala 10:8:@5792.6]
  assign _GEN_57 = _T_2492 % 5'h10; // @[util.scala 10:14:@5793.6]
  assign _T_2493 = _GEN_57[4:0]; // @[util.scala 10:14:@5793.6]
  assign _T_2494 = _T_2493 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5794.6]
  assign _T_2495 = io_storeEmpty & _T_2494; // @[AxiLoadQueue.scala 96:50:@5795.6]
  assign _T_2497 = _T_2495 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5796.6]
  assign _T_2499 = previousStoreHead <= offsetQ_9; // @[AxiLoadQueue.scala 101:36:@5804.8]
  assign _T_2500 = offsetQ_9 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5805.8]
  assign _T_2501 = _T_2499 & _T_2500; // @[AxiLoadQueue.scala 101:61:@5806.8]
  assign _T_2504 = io_storeHead <= offsetQ_9; // @[AxiLoadQueue.scala 103:69:@5812.10]
  assign _T_2505 = offsetQ_9 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5813.10]
  assign _T_2506 = _T_2504 & _T_2505; // @[AxiLoadQueue.scala 103:94:@5814.10]
  assign _T_2508 = _T_2506 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5815.10]
  assign _T_2509 = _T_2233 & _T_2508; // @[AxiLoadQueue.scala 103:51:@5816.10]
  assign _GEN_740 = _T_2509 ? 1'h0 : checkBits_9; // @[AxiLoadQueue.scala 104:53:@5817.10]
  assign _GEN_741 = _T_2501 ? 1'h0 : _GEN_740; // @[AxiLoadQueue.scala 101:102:@5807.8]
  assign _GEN_742 = io_storeEmpty ? 1'h0 : _GEN_741; // @[AxiLoadQueue.scala 99:27:@5800.6]
  assign _GEN_743 = initBits_9 ? _T_2497 : _GEN_742; // @[AxiLoadQueue.scala 95:34:@5785.4]
  assign _T_2522 = _GEN_355 + 4'h1; // @[util.scala 10:8:@5828.6]
  assign _GEN_58 = _T_2522 % 5'h10; // @[util.scala 10:14:@5829.6]
  assign _T_2523 = _GEN_58[4:0]; // @[util.scala 10:14:@5829.6]
  assign _T_2524 = _T_2523 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5830.6]
  assign _T_2525 = io_storeEmpty & _T_2524; // @[AxiLoadQueue.scala 96:50:@5831.6]
  assign _T_2527 = _T_2525 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5832.6]
  assign _T_2529 = previousStoreHead <= offsetQ_10; // @[AxiLoadQueue.scala 101:36:@5840.8]
  assign _T_2530 = offsetQ_10 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5841.8]
  assign _T_2531 = _T_2529 & _T_2530; // @[AxiLoadQueue.scala 101:61:@5842.8]
  assign _T_2534 = io_storeHead <= offsetQ_10; // @[AxiLoadQueue.scala 103:69:@5848.10]
  assign _T_2535 = offsetQ_10 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5849.10]
  assign _T_2536 = _T_2534 & _T_2535; // @[AxiLoadQueue.scala 103:94:@5850.10]
  assign _T_2538 = _T_2536 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5851.10]
  assign _T_2539 = _T_2233 & _T_2538; // @[AxiLoadQueue.scala 103:51:@5852.10]
  assign _GEN_760 = _T_2539 ? 1'h0 : checkBits_10; // @[AxiLoadQueue.scala 104:53:@5853.10]
  assign _GEN_761 = _T_2531 ? 1'h0 : _GEN_760; // @[AxiLoadQueue.scala 101:102:@5843.8]
  assign _GEN_762 = io_storeEmpty ? 1'h0 : _GEN_761; // @[AxiLoadQueue.scala 99:27:@5836.6]
  assign _GEN_763 = initBits_10 ? _T_2527 : _GEN_762; // @[AxiLoadQueue.scala 95:34:@5821.4]
  assign _T_2552 = _GEN_389 + 4'h1; // @[util.scala 10:8:@5864.6]
  assign _GEN_59 = _T_2552 % 5'h10; // @[util.scala 10:14:@5865.6]
  assign _T_2553 = _GEN_59[4:0]; // @[util.scala 10:14:@5865.6]
  assign _T_2554 = _T_2553 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5866.6]
  assign _T_2555 = io_storeEmpty & _T_2554; // @[AxiLoadQueue.scala 96:50:@5867.6]
  assign _T_2557 = _T_2555 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5868.6]
  assign _T_2559 = previousStoreHead <= offsetQ_11; // @[AxiLoadQueue.scala 101:36:@5876.8]
  assign _T_2560 = offsetQ_11 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5877.8]
  assign _T_2561 = _T_2559 & _T_2560; // @[AxiLoadQueue.scala 101:61:@5878.8]
  assign _T_2564 = io_storeHead <= offsetQ_11; // @[AxiLoadQueue.scala 103:69:@5884.10]
  assign _T_2565 = offsetQ_11 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5885.10]
  assign _T_2566 = _T_2564 & _T_2565; // @[AxiLoadQueue.scala 103:94:@5886.10]
  assign _T_2568 = _T_2566 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5887.10]
  assign _T_2569 = _T_2233 & _T_2568; // @[AxiLoadQueue.scala 103:51:@5888.10]
  assign _GEN_780 = _T_2569 ? 1'h0 : checkBits_11; // @[AxiLoadQueue.scala 104:53:@5889.10]
  assign _GEN_781 = _T_2561 ? 1'h0 : _GEN_780; // @[AxiLoadQueue.scala 101:102:@5879.8]
  assign _GEN_782 = io_storeEmpty ? 1'h0 : _GEN_781; // @[AxiLoadQueue.scala 99:27:@5872.6]
  assign _GEN_783 = initBits_11 ? _T_2557 : _GEN_782; // @[AxiLoadQueue.scala 95:34:@5857.4]
  assign _T_2582 = _GEN_423 + 4'h1; // @[util.scala 10:8:@5900.6]
  assign _GEN_60 = _T_2582 % 5'h10; // @[util.scala 10:14:@5901.6]
  assign _T_2583 = _GEN_60[4:0]; // @[util.scala 10:14:@5901.6]
  assign _T_2584 = _T_2583 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5902.6]
  assign _T_2585 = io_storeEmpty & _T_2584; // @[AxiLoadQueue.scala 96:50:@5903.6]
  assign _T_2587 = _T_2585 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5904.6]
  assign _T_2589 = previousStoreHead <= offsetQ_12; // @[AxiLoadQueue.scala 101:36:@5912.8]
  assign _T_2590 = offsetQ_12 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5913.8]
  assign _T_2591 = _T_2589 & _T_2590; // @[AxiLoadQueue.scala 101:61:@5914.8]
  assign _T_2594 = io_storeHead <= offsetQ_12; // @[AxiLoadQueue.scala 103:69:@5920.10]
  assign _T_2595 = offsetQ_12 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5921.10]
  assign _T_2596 = _T_2594 & _T_2595; // @[AxiLoadQueue.scala 103:94:@5922.10]
  assign _T_2598 = _T_2596 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5923.10]
  assign _T_2599 = _T_2233 & _T_2598; // @[AxiLoadQueue.scala 103:51:@5924.10]
  assign _GEN_800 = _T_2599 ? 1'h0 : checkBits_12; // @[AxiLoadQueue.scala 104:53:@5925.10]
  assign _GEN_801 = _T_2591 ? 1'h0 : _GEN_800; // @[AxiLoadQueue.scala 101:102:@5915.8]
  assign _GEN_802 = io_storeEmpty ? 1'h0 : _GEN_801; // @[AxiLoadQueue.scala 99:27:@5908.6]
  assign _GEN_803 = initBits_12 ? _T_2587 : _GEN_802; // @[AxiLoadQueue.scala 95:34:@5893.4]
  assign _T_2612 = _GEN_457 + 4'h1; // @[util.scala 10:8:@5936.6]
  assign _GEN_61 = _T_2612 % 5'h10; // @[util.scala 10:14:@5937.6]
  assign _T_2613 = _GEN_61[4:0]; // @[util.scala 10:14:@5937.6]
  assign _T_2614 = _T_2613 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5938.6]
  assign _T_2615 = io_storeEmpty & _T_2614; // @[AxiLoadQueue.scala 96:50:@5939.6]
  assign _T_2617 = _T_2615 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5940.6]
  assign _T_2619 = previousStoreHead <= offsetQ_13; // @[AxiLoadQueue.scala 101:36:@5948.8]
  assign _T_2620 = offsetQ_13 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5949.8]
  assign _T_2621 = _T_2619 & _T_2620; // @[AxiLoadQueue.scala 101:61:@5950.8]
  assign _T_2624 = io_storeHead <= offsetQ_13; // @[AxiLoadQueue.scala 103:69:@5956.10]
  assign _T_2625 = offsetQ_13 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5957.10]
  assign _T_2626 = _T_2624 & _T_2625; // @[AxiLoadQueue.scala 103:94:@5958.10]
  assign _T_2628 = _T_2626 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5959.10]
  assign _T_2629 = _T_2233 & _T_2628; // @[AxiLoadQueue.scala 103:51:@5960.10]
  assign _GEN_820 = _T_2629 ? 1'h0 : checkBits_13; // @[AxiLoadQueue.scala 104:53:@5961.10]
  assign _GEN_821 = _T_2621 ? 1'h0 : _GEN_820; // @[AxiLoadQueue.scala 101:102:@5951.8]
  assign _GEN_822 = io_storeEmpty ? 1'h0 : _GEN_821; // @[AxiLoadQueue.scala 99:27:@5944.6]
  assign _GEN_823 = initBits_13 ? _T_2617 : _GEN_822; // @[AxiLoadQueue.scala 95:34:@5929.4]
  assign _T_2642 = _GEN_491 + 4'h1; // @[util.scala 10:8:@5972.6]
  assign _GEN_62 = _T_2642 % 5'h10; // @[util.scala 10:14:@5973.6]
  assign _T_2643 = _GEN_62[4:0]; // @[util.scala 10:14:@5973.6]
  assign _T_2644 = _T_2643 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@5974.6]
  assign _T_2645 = io_storeEmpty & _T_2644; // @[AxiLoadQueue.scala 96:50:@5975.6]
  assign _T_2647 = _T_2645 == 1'h0; // @[AxiLoadQueue.scala 96:34:@5976.6]
  assign _T_2649 = previousStoreHead <= offsetQ_14; // @[AxiLoadQueue.scala 101:36:@5984.8]
  assign _T_2650 = offsetQ_14 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@5985.8]
  assign _T_2651 = _T_2649 & _T_2650; // @[AxiLoadQueue.scala 101:61:@5986.8]
  assign _T_2654 = io_storeHead <= offsetQ_14; // @[AxiLoadQueue.scala 103:69:@5992.10]
  assign _T_2655 = offsetQ_14 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@5993.10]
  assign _T_2656 = _T_2654 & _T_2655; // @[AxiLoadQueue.scala 103:94:@5994.10]
  assign _T_2658 = _T_2656 == 1'h0; // @[AxiLoadQueue.scala 103:54:@5995.10]
  assign _T_2659 = _T_2233 & _T_2658; // @[AxiLoadQueue.scala 103:51:@5996.10]
  assign _GEN_840 = _T_2659 ? 1'h0 : checkBits_14; // @[AxiLoadQueue.scala 104:53:@5997.10]
  assign _GEN_841 = _T_2651 ? 1'h0 : _GEN_840; // @[AxiLoadQueue.scala 101:102:@5987.8]
  assign _GEN_842 = io_storeEmpty ? 1'h0 : _GEN_841; // @[AxiLoadQueue.scala 99:27:@5980.6]
  assign _GEN_843 = initBits_14 ? _T_2647 : _GEN_842; // @[AxiLoadQueue.scala 95:34:@5965.4]
  assign _T_2672 = _GEN_525 + 4'h1; // @[util.scala 10:8:@6008.6]
  assign _GEN_63 = _T_2672 % 5'h10; // @[util.scala 10:14:@6009.6]
  assign _T_2673 = _GEN_63[4:0]; // @[util.scala 10:14:@6009.6]
  assign _T_2674 = _T_2673 == _GEN_2341; // @[AxiLoadQueue.scala 97:56:@6010.6]
  assign _T_2675 = io_storeEmpty & _T_2674; // @[AxiLoadQueue.scala 96:50:@6011.6]
  assign _T_2677 = _T_2675 == 1'h0; // @[AxiLoadQueue.scala 96:34:@6012.6]
  assign _T_2679 = previousStoreHead <= offsetQ_15; // @[AxiLoadQueue.scala 101:36:@6020.8]
  assign _T_2680 = offsetQ_15 < io_storeHead; // @[AxiLoadQueue.scala 101:86:@6021.8]
  assign _T_2681 = _T_2679 & _T_2680; // @[AxiLoadQueue.scala 101:61:@6022.8]
  assign _T_2684 = io_storeHead <= offsetQ_15; // @[AxiLoadQueue.scala 103:69:@6028.10]
  assign _T_2685 = offsetQ_15 < previousStoreHead; // @[AxiLoadQueue.scala 104:31:@6029.10]
  assign _T_2686 = _T_2684 & _T_2685; // @[AxiLoadQueue.scala 103:94:@6030.10]
  assign _T_2688 = _T_2686 == 1'h0; // @[AxiLoadQueue.scala 103:54:@6031.10]
  assign _T_2689 = _T_2233 & _T_2688; // @[AxiLoadQueue.scala 103:51:@6032.10]
  assign _GEN_860 = _T_2689 ? 1'h0 : checkBits_15; // @[AxiLoadQueue.scala 104:53:@6033.10]
  assign _GEN_861 = _T_2681 ? 1'h0 : _GEN_860; // @[AxiLoadQueue.scala 101:102:@6023.8]
  assign _GEN_862 = io_storeEmpty ? 1'h0 : _GEN_861; // @[AxiLoadQueue.scala 99:27:@6016.6]
  assign _GEN_863 = initBits_15 ? _T_2677 : _GEN_862; // @[AxiLoadQueue.scala 95:34:@6001.4]
  assign _T_2693 = 16'h1 << io_storeHead; // @[OneHot.scala 52:12:@6038.4]
  assign _T_2695 = _T_2693[0]; // @[util.scala 60:60:@6040.4]
  assign _T_2696 = _T_2693[1]; // @[util.scala 60:60:@6041.4]
  assign _T_2697 = _T_2693[2]; // @[util.scala 60:60:@6042.4]
  assign _T_2698 = _T_2693[3]; // @[util.scala 60:60:@6043.4]
  assign _T_2699 = _T_2693[4]; // @[util.scala 60:60:@6044.4]
  assign _T_2700 = _T_2693[5]; // @[util.scala 60:60:@6045.4]
  assign _T_2701 = _T_2693[6]; // @[util.scala 60:60:@6046.4]
  assign _T_2702 = _T_2693[7]; // @[util.scala 60:60:@6047.4]
  assign _T_2703 = _T_2693[8]; // @[util.scala 60:60:@6048.4]
  assign _T_2704 = _T_2693[9]; // @[util.scala 60:60:@6049.4]
  assign _T_2705 = _T_2693[10]; // @[util.scala 60:60:@6050.4]
  assign _T_2706 = _T_2693[11]; // @[util.scala 60:60:@6051.4]
  assign _T_2707 = _T_2693[12]; // @[util.scala 60:60:@6052.4]
  assign _T_2708 = _T_2693[13]; // @[util.scala 60:60:@6053.4]
  assign _T_2709 = _T_2693[14]; // @[util.scala 60:60:@6054.4]
  assign _T_2710 = _T_2693[15]; // @[util.scala 60:60:@6055.4]
  assign _T_4841 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0}; // @[Mux.scala 19:72:@7579.4]
  assign _T_4848 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8}; // @[Mux.scala 19:72:@7586.4]
  assign _T_4849 = {io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,_T_4841}; // @[Mux.scala 19:72:@7587.4]
  assign _T_4851 = _T_2695 ? _T_4849 : 512'h0; // @[Mux.scala 19:72:@7588.4]
  assign _T_4858 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1}; // @[Mux.scala 19:72:@7595.4]
  assign _T_4865 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9}; // @[Mux.scala 19:72:@7602.4]
  assign _T_4866 = {io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,_T_4858}; // @[Mux.scala 19:72:@7603.4]
  assign _T_4868 = _T_2696 ? _T_4866 : 512'h0; // @[Mux.scala 19:72:@7604.4]
  assign _T_4875 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2}; // @[Mux.scala 19:72:@7611.4]
  assign _T_4882 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10}; // @[Mux.scala 19:72:@7618.4]
  assign _T_4883 = {io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,_T_4875}; // @[Mux.scala 19:72:@7619.4]
  assign _T_4885 = _T_2697 ? _T_4883 : 512'h0; // @[Mux.scala 19:72:@7620.4]
  assign _T_4892 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3}; // @[Mux.scala 19:72:@7627.4]
  assign _T_4899 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11}; // @[Mux.scala 19:72:@7634.4]
  assign _T_4900 = {io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,_T_4892}; // @[Mux.scala 19:72:@7635.4]
  assign _T_4902 = _T_2698 ? _T_4900 : 512'h0; // @[Mux.scala 19:72:@7636.4]
  assign _T_4909 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4}; // @[Mux.scala 19:72:@7643.4]
  assign _T_4916 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12}; // @[Mux.scala 19:72:@7650.4]
  assign _T_4917 = {io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,_T_4909}; // @[Mux.scala 19:72:@7651.4]
  assign _T_4919 = _T_2699 ? _T_4917 : 512'h0; // @[Mux.scala 19:72:@7652.4]
  assign _T_4926 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5}; // @[Mux.scala 19:72:@7659.4]
  assign _T_4933 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13}; // @[Mux.scala 19:72:@7666.4]
  assign _T_4934 = {io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,io_storeDataQueue_13,_T_4926}; // @[Mux.scala 19:72:@7667.4]
  assign _T_4936 = _T_2700 ? _T_4934 : 512'h0; // @[Mux.scala 19:72:@7668.4]
  assign _T_4943 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6}; // @[Mux.scala 19:72:@7675.4]
  assign _T_4950 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14}; // @[Mux.scala 19:72:@7682.4]
  assign _T_4951 = {io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,io_storeDataQueue_14,_T_4943}; // @[Mux.scala 19:72:@7683.4]
  assign _T_4953 = _T_2701 ? _T_4951 : 512'h0; // @[Mux.scala 19:72:@7684.4]
  assign _T_4960 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7}; // @[Mux.scala 19:72:@7691.4]
  assign _T_4967 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15}; // @[Mux.scala 19:72:@7698.4]
  assign _T_4968 = {io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,io_storeDataQueue_15,_T_4960}; // @[Mux.scala 19:72:@7699.4]
  assign _T_4970 = _T_2702 ? _T_4968 : 512'h0; // @[Mux.scala 19:72:@7700.4]
  assign _T_4985 = {io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,io_storeDataQueue_0,_T_4848}; // @[Mux.scala 19:72:@7715.4]
  assign _T_4987 = _T_2703 ? _T_4985 : 512'h0; // @[Mux.scala 19:72:@7716.4]
  assign _T_5002 = {io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,io_storeDataQueue_1,_T_4865}; // @[Mux.scala 19:72:@7731.4]
  assign _T_5004 = _T_2704 ? _T_5002 : 512'h0; // @[Mux.scala 19:72:@7732.4]
  assign _T_5019 = {io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,io_storeDataQueue_2,_T_4882}; // @[Mux.scala 19:72:@7747.4]
  assign _T_5021 = _T_2705 ? _T_5019 : 512'h0; // @[Mux.scala 19:72:@7748.4]
  assign _T_5036 = {io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,io_storeDataQueue_3,_T_4899}; // @[Mux.scala 19:72:@7763.4]
  assign _T_5038 = _T_2706 ? _T_5036 : 512'h0; // @[Mux.scala 19:72:@7764.4]
  assign _T_5053 = {io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,io_storeDataQueue_4,_T_4916}; // @[Mux.scala 19:72:@7779.4]
  assign _T_5055 = _T_2707 ? _T_5053 : 512'h0; // @[Mux.scala 19:72:@7780.4]
  assign _T_5070 = {io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,io_storeDataQueue_5,_T_4933}; // @[Mux.scala 19:72:@7795.4]
  assign _T_5072 = _T_2708 ? _T_5070 : 512'h0; // @[Mux.scala 19:72:@7796.4]
  assign _T_5087 = {io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,io_storeDataQueue_6,_T_4950}; // @[Mux.scala 19:72:@7811.4]
  assign _T_5089 = _T_2709 ? _T_5087 : 512'h0; // @[Mux.scala 19:72:@7812.4]
  assign _T_5104 = {io_storeDataQueue_14,io_storeDataQueue_13,io_storeDataQueue_12,io_storeDataQueue_11,io_storeDataQueue_10,io_storeDataQueue_9,io_storeDataQueue_8,io_storeDataQueue_7,_T_4967}; // @[Mux.scala 19:72:@7827.4]
  assign _T_5106 = _T_2710 ? _T_5104 : 512'h0; // @[Mux.scala 19:72:@7828.4]
  assign _T_5107 = _T_4851 | _T_4868; // @[Mux.scala 19:72:@7829.4]
  assign _T_5108 = _T_5107 | _T_4885; // @[Mux.scala 19:72:@7830.4]
  assign _T_5109 = _T_5108 | _T_4902; // @[Mux.scala 19:72:@7831.4]
  assign _T_5110 = _T_5109 | _T_4919; // @[Mux.scala 19:72:@7832.4]
  assign _T_5111 = _T_5110 | _T_4936; // @[Mux.scala 19:72:@7833.4]
  assign _T_5112 = _T_5111 | _T_4953; // @[Mux.scala 19:72:@7834.4]
  assign _T_5113 = _T_5112 | _T_4970; // @[Mux.scala 19:72:@7835.4]
  assign _T_5114 = _T_5113 | _T_4987; // @[Mux.scala 19:72:@7836.4]
  assign _T_5115 = _T_5114 | _T_5004; // @[Mux.scala 19:72:@7837.4]
  assign _T_5116 = _T_5115 | _T_5021; // @[Mux.scala 19:72:@7838.4]
  assign _T_5117 = _T_5116 | _T_5038; // @[Mux.scala 19:72:@7839.4]
  assign _T_5118 = _T_5117 | _T_5055; // @[Mux.scala 19:72:@7840.4]
  assign _T_5119 = _T_5118 | _T_5072; // @[Mux.scala 19:72:@7841.4]
  assign _T_5120 = _T_5119 | _T_5089; // @[Mux.scala 19:72:@7842.4]
  assign _T_5121 = _T_5120 | _T_5106; // @[Mux.scala 19:72:@7843.4]
  assign _T_5698 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0}; // @[Mux.scala 19:72:@8193.4]
  assign _T_5705 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8}; // @[Mux.scala 19:72:@8200.4]
  assign _T_5706 = {io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,_T_5698}; // @[Mux.scala 19:72:@8201.4]
  assign _T_5708 = _T_2695 ? _T_5706 : 16'h0; // @[Mux.scala 19:72:@8202.4]
  assign _T_5715 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1}; // @[Mux.scala 19:72:@8209.4]
  assign _T_5722 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9}; // @[Mux.scala 19:72:@8216.4]
  assign _T_5723 = {io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,_T_5715}; // @[Mux.scala 19:72:@8217.4]
  assign _T_5725 = _T_2696 ? _T_5723 : 16'h0; // @[Mux.scala 19:72:@8218.4]
  assign _T_5732 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2}; // @[Mux.scala 19:72:@8225.4]
  assign _T_5739 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10}; // @[Mux.scala 19:72:@8232.4]
  assign _T_5740 = {io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,_T_5732}; // @[Mux.scala 19:72:@8233.4]
  assign _T_5742 = _T_2697 ? _T_5740 : 16'h0; // @[Mux.scala 19:72:@8234.4]
  assign _T_5749 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3}; // @[Mux.scala 19:72:@8241.4]
  assign _T_5756 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11}; // @[Mux.scala 19:72:@8248.4]
  assign _T_5757 = {io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,_T_5749}; // @[Mux.scala 19:72:@8249.4]
  assign _T_5759 = _T_2698 ? _T_5757 : 16'h0; // @[Mux.scala 19:72:@8250.4]
  assign _T_5766 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4}; // @[Mux.scala 19:72:@8257.4]
  assign _T_5773 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12}; // @[Mux.scala 19:72:@8264.4]
  assign _T_5774 = {io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,_T_5766}; // @[Mux.scala 19:72:@8265.4]
  assign _T_5776 = _T_2699 ? _T_5774 : 16'h0; // @[Mux.scala 19:72:@8266.4]
  assign _T_5783 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5}; // @[Mux.scala 19:72:@8273.4]
  assign _T_5790 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13}; // @[Mux.scala 19:72:@8280.4]
  assign _T_5791 = {io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,io_storeDataDone_13,_T_5783}; // @[Mux.scala 19:72:@8281.4]
  assign _T_5793 = _T_2700 ? _T_5791 : 16'h0; // @[Mux.scala 19:72:@8282.4]
  assign _T_5800 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6}; // @[Mux.scala 19:72:@8289.4]
  assign _T_5807 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14}; // @[Mux.scala 19:72:@8296.4]
  assign _T_5808 = {io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,io_storeDataDone_14,_T_5800}; // @[Mux.scala 19:72:@8297.4]
  assign _T_5810 = _T_2701 ? _T_5808 : 16'h0; // @[Mux.scala 19:72:@8298.4]
  assign _T_5817 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7}; // @[Mux.scala 19:72:@8305.4]
  assign _T_5824 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15}; // @[Mux.scala 19:72:@8312.4]
  assign _T_5825 = {io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,io_storeDataDone_15,_T_5817}; // @[Mux.scala 19:72:@8313.4]
  assign _T_5827 = _T_2702 ? _T_5825 : 16'h0; // @[Mux.scala 19:72:@8314.4]
  assign _T_5842 = {io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,io_storeDataDone_0,_T_5705}; // @[Mux.scala 19:72:@8329.4]
  assign _T_5844 = _T_2703 ? _T_5842 : 16'h0; // @[Mux.scala 19:72:@8330.4]
  assign _T_5859 = {io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,io_storeDataDone_1,_T_5722}; // @[Mux.scala 19:72:@8345.4]
  assign _T_5861 = _T_2704 ? _T_5859 : 16'h0; // @[Mux.scala 19:72:@8346.4]
  assign _T_5876 = {io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,io_storeDataDone_2,_T_5739}; // @[Mux.scala 19:72:@8361.4]
  assign _T_5878 = _T_2705 ? _T_5876 : 16'h0; // @[Mux.scala 19:72:@8362.4]
  assign _T_5893 = {io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,io_storeDataDone_3,_T_5756}; // @[Mux.scala 19:72:@8377.4]
  assign _T_5895 = _T_2706 ? _T_5893 : 16'h0; // @[Mux.scala 19:72:@8378.4]
  assign _T_5910 = {io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,io_storeDataDone_4,_T_5773}; // @[Mux.scala 19:72:@8393.4]
  assign _T_5912 = _T_2707 ? _T_5910 : 16'h0; // @[Mux.scala 19:72:@8394.4]
  assign _T_5927 = {io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,io_storeDataDone_5,_T_5790}; // @[Mux.scala 19:72:@8409.4]
  assign _T_5929 = _T_2708 ? _T_5927 : 16'h0; // @[Mux.scala 19:72:@8410.4]
  assign _T_5944 = {io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,io_storeDataDone_6,_T_5807}; // @[Mux.scala 19:72:@8425.4]
  assign _T_5946 = _T_2709 ? _T_5944 : 16'h0; // @[Mux.scala 19:72:@8426.4]
  assign _T_5961 = {io_storeDataDone_14,io_storeDataDone_13,io_storeDataDone_12,io_storeDataDone_11,io_storeDataDone_10,io_storeDataDone_9,io_storeDataDone_8,io_storeDataDone_7,_T_5824}; // @[Mux.scala 19:72:@8441.4]
  assign _T_5963 = _T_2710 ? _T_5961 : 16'h0; // @[Mux.scala 19:72:@8442.4]
  assign _T_5964 = _T_5708 | _T_5725; // @[Mux.scala 19:72:@8443.4]
  assign _T_5965 = _T_5964 | _T_5742; // @[Mux.scala 19:72:@8444.4]
  assign _T_5966 = _T_5965 | _T_5759; // @[Mux.scala 19:72:@8445.4]
  assign _T_5967 = _T_5966 | _T_5776; // @[Mux.scala 19:72:@8446.4]
  assign _T_5968 = _T_5967 | _T_5793; // @[Mux.scala 19:72:@8447.4]
  assign _T_5969 = _T_5968 | _T_5810; // @[Mux.scala 19:72:@8448.4]
  assign _T_5970 = _T_5969 | _T_5827; // @[Mux.scala 19:72:@8449.4]
  assign _T_5971 = _T_5970 | _T_5844; // @[Mux.scala 19:72:@8450.4]
  assign _T_5972 = _T_5971 | _T_5861; // @[Mux.scala 19:72:@8451.4]
  assign _T_5973 = _T_5972 | _T_5878; // @[Mux.scala 19:72:@8452.4]
  assign _T_5974 = _T_5973 | _T_5895; // @[Mux.scala 19:72:@8453.4]
  assign _T_5975 = _T_5974 | _T_5912; // @[Mux.scala 19:72:@8454.4]
  assign _T_5976 = _T_5975 | _T_5929; // @[Mux.scala 19:72:@8455.4]
  assign _T_5977 = _T_5976 | _T_5946; // @[Mux.scala 19:72:@8456.4]
  assign _T_5978 = _T_5977 | _T_5963; // @[Mux.scala 19:72:@8457.4]
  assign _T_6119 = io_storeHead < io_storeTail; // @[AxiLoadQueue.scala 121:105:@8493.4]
  assign _T_6121 = io_storeHead <= 4'h0; // @[AxiLoadQueue.scala 122:18:@8494.4]
  assign _T_6123 = 4'h0 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8495.4]
  assign _T_6124 = _T_6121 & _T_6123; // @[AxiLoadQueue.scala 122:27:@8496.4]
  assign _T_6126 = io_storeEmpty == 1'h0; // @[AxiLoadQueue.scala 122:52:@8497.4]
  assign _T_6128 = io_storeTail <= 4'h0; // @[AxiLoadQueue.scala 122:85:@8498.4]
  assign _T_6130 = 4'h0 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8499.4]
  assign _T_6131 = _T_6128 & _T_6130; // @[AxiLoadQueue.scala 122:94:@8500.4]
  assign _T_6133 = _T_6131 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8501.4]
  assign _T_6134 = _T_6126 & _T_6133; // @[AxiLoadQueue.scala 122:67:@8502.4]
  assign validEntriesInStoreQ_0 = _T_6119 ? _T_6124 : _T_6134; // @[AxiLoadQueue.scala 121:91:@8503.4]
  assign _T_6138 = io_storeHead <= 4'h1; // @[AxiLoadQueue.scala 122:18:@8505.4]
  assign _T_6140 = 4'h1 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8506.4]
  assign _T_6141 = _T_6138 & _T_6140; // @[AxiLoadQueue.scala 122:27:@8507.4]
  assign _T_6145 = io_storeTail <= 4'h1; // @[AxiLoadQueue.scala 122:85:@8509.4]
  assign _T_6147 = 4'h1 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8510.4]
  assign _T_6148 = _T_6145 & _T_6147; // @[AxiLoadQueue.scala 122:94:@8511.4]
  assign _T_6150 = _T_6148 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8512.4]
  assign _T_6151 = _T_6126 & _T_6150; // @[AxiLoadQueue.scala 122:67:@8513.4]
  assign validEntriesInStoreQ_1 = _T_6119 ? _T_6141 : _T_6151; // @[AxiLoadQueue.scala 121:91:@8514.4]
  assign _T_6155 = io_storeHead <= 4'h2; // @[AxiLoadQueue.scala 122:18:@8516.4]
  assign _T_6157 = 4'h2 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8517.4]
  assign _T_6158 = _T_6155 & _T_6157; // @[AxiLoadQueue.scala 122:27:@8518.4]
  assign _T_6162 = io_storeTail <= 4'h2; // @[AxiLoadQueue.scala 122:85:@8520.4]
  assign _T_6164 = 4'h2 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8521.4]
  assign _T_6165 = _T_6162 & _T_6164; // @[AxiLoadQueue.scala 122:94:@8522.4]
  assign _T_6167 = _T_6165 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8523.4]
  assign _T_6168 = _T_6126 & _T_6167; // @[AxiLoadQueue.scala 122:67:@8524.4]
  assign validEntriesInStoreQ_2 = _T_6119 ? _T_6158 : _T_6168; // @[AxiLoadQueue.scala 121:91:@8525.4]
  assign _T_6172 = io_storeHead <= 4'h3; // @[AxiLoadQueue.scala 122:18:@8527.4]
  assign _T_6174 = 4'h3 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8528.4]
  assign _T_6175 = _T_6172 & _T_6174; // @[AxiLoadQueue.scala 122:27:@8529.4]
  assign _T_6179 = io_storeTail <= 4'h3; // @[AxiLoadQueue.scala 122:85:@8531.4]
  assign _T_6181 = 4'h3 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8532.4]
  assign _T_6182 = _T_6179 & _T_6181; // @[AxiLoadQueue.scala 122:94:@8533.4]
  assign _T_6184 = _T_6182 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8534.4]
  assign _T_6185 = _T_6126 & _T_6184; // @[AxiLoadQueue.scala 122:67:@8535.4]
  assign validEntriesInStoreQ_3 = _T_6119 ? _T_6175 : _T_6185; // @[AxiLoadQueue.scala 121:91:@8536.4]
  assign _T_6189 = io_storeHead <= 4'h4; // @[AxiLoadQueue.scala 122:18:@8538.4]
  assign _T_6191 = 4'h4 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8539.4]
  assign _T_6192 = _T_6189 & _T_6191; // @[AxiLoadQueue.scala 122:27:@8540.4]
  assign _T_6196 = io_storeTail <= 4'h4; // @[AxiLoadQueue.scala 122:85:@8542.4]
  assign _T_6198 = 4'h4 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8543.4]
  assign _T_6199 = _T_6196 & _T_6198; // @[AxiLoadQueue.scala 122:94:@8544.4]
  assign _T_6201 = _T_6199 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8545.4]
  assign _T_6202 = _T_6126 & _T_6201; // @[AxiLoadQueue.scala 122:67:@8546.4]
  assign validEntriesInStoreQ_4 = _T_6119 ? _T_6192 : _T_6202; // @[AxiLoadQueue.scala 121:91:@8547.4]
  assign _T_6206 = io_storeHead <= 4'h5; // @[AxiLoadQueue.scala 122:18:@8549.4]
  assign _T_6208 = 4'h5 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8550.4]
  assign _T_6209 = _T_6206 & _T_6208; // @[AxiLoadQueue.scala 122:27:@8551.4]
  assign _T_6213 = io_storeTail <= 4'h5; // @[AxiLoadQueue.scala 122:85:@8553.4]
  assign _T_6215 = 4'h5 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8554.4]
  assign _T_6216 = _T_6213 & _T_6215; // @[AxiLoadQueue.scala 122:94:@8555.4]
  assign _T_6218 = _T_6216 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8556.4]
  assign _T_6219 = _T_6126 & _T_6218; // @[AxiLoadQueue.scala 122:67:@8557.4]
  assign validEntriesInStoreQ_5 = _T_6119 ? _T_6209 : _T_6219; // @[AxiLoadQueue.scala 121:91:@8558.4]
  assign _T_6223 = io_storeHead <= 4'h6; // @[AxiLoadQueue.scala 122:18:@8560.4]
  assign _T_6225 = 4'h6 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8561.4]
  assign _T_6226 = _T_6223 & _T_6225; // @[AxiLoadQueue.scala 122:27:@8562.4]
  assign _T_6230 = io_storeTail <= 4'h6; // @[AxiLoadQueue.scala 122:85:@8564.4]
  assign _T_6232 = 4'h6 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8565.4]
  assign _T_6233 = _T_6230 & _T_6232; // @[AxiLoadQueue.scala 122:94:@8566.4]
  assign _T_6235 = _T_6233 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8567.4]
  assign _T_6236 = _T_6126 & _T_6235; // @[AxiLoadQueue.scala 122:67:@8568.4]
  assign validEntriesInStoreQ_6 = _T_6119 ? _T_6226 : _T_6236; // @[AxiLoadQueue.scala 121:91:@8569.4]
  assign _T_6240 = io_storeHead <= 4'h7; // @[AxiLoadQueue.scala 122:18:@8571.4]
  assign _T_6242 = 4'h7 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8572.4]
  assign _T_6243 = _T_6240 & _T_6242; // @[AxiLoadQueue.scala 122:27:@8573.4]
  assign _T_6247 = io_storeTail <= 4'h7; // @[AxiLoadQueue.scala 122:85:@8575.4]
  assign _T_6249 = 4'h7 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8576.4]
  assign _T_6250 = _T_6247 & _T_6249; // @[AxiLoadQueue.scala 122:94:@8577.4]
  assign _T_6252 = _T_6250 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8578.4]
  assign _T_6253 = _T_6126 & _T_6252; // @[AxiLoadQueue.scala 122:67:@8579.4]
  assign validEntriesInStoreQ_7 = _T_6119 ? _T_6243 : _T_6253; // @[AxiLoadQueue.scala 121:91:@8580.4]
  assign _T_6257 = io_storeHead <= 4'h8; // @[AxiLoadQueue.scala 122:18:@8582.4]
  assign _T_6259 = 4'h8 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8583.4]
  assign _T_6260 = _T_6257 & _T_6259; // @[AxiLoadQueue.scala 122:27:@8584.4]
  assign _T_6264 = io_storeTail <= 4'h8; // @[AxiLoadQueue.scala 122:85:@8586.4]
  assign _T_6266 = 4'h8 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8587.4]
  assign _T_6267 = _T_6264 & _T_6266; // @[AxiLoadQueue.scala 122:94:@8588.4]
  assign _T_6269 = _T_6267 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8589.4]
  assign _T_6270 = _T_6126 & _T_6269; // @[AxiLoadQueue.scala 122:67:@8590.4]
  assign validEntriesInStoreQ_8 = _T_6119 ? _T_6260 : _T_6270; // @[AxiLoadQueue.scala 121:91:@8591.4]
  assign _T_6274 = io_storeHead <= 4'h9; // @[AxiLoadQueue.scala 122:18:@8593.4]
  assign _T_6276 = 4'h9 < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8594.4]
  assign _T_6277 = _T_6274 & _T_6276; // @[AxiLoadQueue.scala 122:27:@8595.4]
  assign _T_6281 = io_storeTail <= 4'h9; // @[AxiLoadQueue.scala 122:85:@8597.4]
  assign _T_6283 = 4'h9 < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8598.4]
  assign _T_6284 = _T_6281 & _T_6283; // @[AxiLoadQueue.scala 122:94:@8599.4]
  assign _T_6286 = _T_6284 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8600.4]
  assign _T_6287 = _T_6126 & _T_6286; // @[AxiLoadQueue.scala 122:67:@8601.4]
  assign validEntriesInStoreQ_9 = _T_6119 ? _T_6277 : _T_6287; // @[AxiLoadQueue.scala 121:91:@8602.4]
  assign _T_6291 = io_storeHead <= 4'ha; // @[AxiLoadQueue.scala 122:18:@8604.4]
  assign _T_6293 = 4'ha < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8605.4]
  assign _T_6294 = _T_6291 & _T_6293; // @[AxiLoadQueue.scala 122:27:@8606.4]
  assign _T_6298 = io_storeTail <= 4'ha; // @[AxiLoadQueue.scala 122:85:@8608.4]
  assign _T_6300 = 4'ha < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8609.4]
  assign _T_6301 = _T_6298 & _T_6300; // @[AxiLoadQueue.scala 122:94:@8610.4]
  assign _T_6303 = _T_6301 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8611.4]
  assign _T_6304 = _T_6126 & _T_6303; // @[AxiLoadQueue.scala 122:67:@8612.4]
  assign validEntriesInStoreQ_10 = _T_6119 ? _T_6294 : _T_6304; // @[AxiLoadQueue.scala 121:91:@8613.4]
  assign _T_6308 = io_storeHead <= 4'hb; // @[AxiLoadQueue.scala 122:18:@8615.4]
  assign _T_6310 = 4'hb < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8616.4]
  assign _T_6311 = _T_6308 & _T_6310; // @[AxiLoadQueue.scala 122:27:@8617.4]
  assign _T_6315 = io_storeTail <= 4'hb; // @[AxiLoadQueue.scala 122:85:@8619.4]
  assign _T_6317 = 4'hb < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8620.4]
  assign _T_6318 = _T_6315 & _T_6317; // @[AxiLoadQueue.scala 122:94:@8621.4]
  assign _T_6320 = _T_6318 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8622.4]
  assign _T_6321 = _T_6126 & _T_6320; // @[AxiLoadQueue.scala 122:67:@8623.4]
  assign validEntriesInStoreQ_11 = _T_6119 ? _T_6311 : _T_6321; // @[AxiLoadQueue.scala 121:91:@8624.4]
  assign _T_6325 = io_storeHead <= 4'hc; // @[AxiLoadQueue.scala 122:18:@8626.4]
  assign _T_6327 = 4'hc < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8627.4]
  assign _T_6328 = _T_6325 & _T_6327; // @[AxiLoadQueue.scala 122:27:@8628.4]
  assign _T_6332 = io_storeTail <= 4'hc; // @[AxiLoadQueue.scala 122:85:@8630.4]
  assign _T_6334 = 4'hc < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8631.4]
  assign _T_6335 = _T_6332 & _T_6334; // @[AxiLoadQueue.scala 122:94:@8632.4]
  assign _T_6337 = _T_6335 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8633.4]
  assign _T_6338 = _T_6126 & _T_6337; // @[AxiLoadQueue.scala 122:67:@8634.4]
  assign validEntriesInStoreQ_12 = _T_6119 ? _T_6328 : _T_6338; // @[AxiLoadQueue.scala 121:91:@8635.4]
  assign _T_6342 = io_storeHead <= 4'hd; // @[AxiLoadQueue.scala 122:18:@8637.4]
  assign _T_6344 = 4'hd < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8638.4]
  assign _T_6345 = _T_6342 & _T_6344; // @[AxiLoadQueue.scala 122:27:@8639.4]
  assign _T_6349 = io_storeTail <= 4'hd; // @[AxiLoadQueue.scala 122:85:@8641.4]
  assign _T_6351 = 4'hd < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8642.4]
  assign _T_6352 = _T_6349 & _T_6351; // @[AxiLoadQueue.scala 122:94:@8643.4]
  assign _T_6354 = _T_6352 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8644.4]
  assign _T_6355 = _T_6126 & _T_6354; // @[AxiLoadQueue.scala 122:67:@8645.4]
  assign validEntriesInStoreQ_13 = _T_6119 ? _T_6345 : _T_6355; // @[AxiLoadQueue.scala 121:91:@8646.4]
  assign _T_6359 = io_storeHead <= 4'he; // @[AxiLoadQueue.scala 122:18:@8648.4]
  assign _T_6361 = 4'he < io_storeTail; // @[AxiLoadQueue.scala 122:36:@8649.4]
  assign _T_6362 = _T_6359 & _T_6361; // @[AxiLoadQueue.scala 122:27:@8650.4]
  assign _T_6366 = io_storeTail <= 4'he; // @[AxiLoadQueue.scala 122:85:@8652.4]
  assign _T_6368 = 4'he < io_storeHead; // @[AxiLoadQueue.scala 122:103:@8653.4]
  assign _T_6369 = _T_6366 & _T_6368; // @[AxiLoadQueue.scala 122:94:@8654.4]
  assign _T_6371 = _T_6369 == 1'h0; // @[AxiLoadQueue.scala 122:70:@8655.4]
  assign _T_6372 = _T_6126 & _T_6371; // @[AxiLoadQueue.scala 122:67:@8656.4]
  assign validEntriesInStoreQ_14 = _T_6119 ? _T_6362 : _T_6372; // @[AxiLoadQueue.scala 121:91:@8657.4]
  assign validEntriesInStoreQ_15 = _T_6119 ? 1'h0 : _T_6126; // @[AxiLoadQueue.scala 121:91:@8668.4]
  assign storesToCheck_0_0 = _T_2234 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@8695.4]
  assign _T_7660 = 4'h1 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8698.4]
  assign _T_7661 = _T_6138 & _T_7660; // @[AxiLoadQueue.scala 130:72:@8699.4]
  assign _T_7663 = offsetQ_0 < 4'h1; // @[AxiLoadQueue.scala 131:33:@8700.4]
  assign _T_7666 = _T_7663 & _T_6147; // @[AxiLoadQueue.scala 131:41:@8702.4]
  assign _T_7668 = _T_7666 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8703.4]
  assign storesToCheck_0_1 = _T_2234 ? _T_7661 : _T_7668; // @[AxiLoadQueue.scala 130:10:@8704.4]
  assign _T_7674 = 4'h2 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8707.4]
  assign _T_7675 = _T_6155 & _T_7674; // @[AxiLoadQueue.scala 130:72:@8708.4]
  assign _T_7677 = offsetQ_0 < 4'h2; // @[AxiLoadQueue.scala 131:33:@8709.4]
  assign _T_7680 = _T_7677 & _T_6164; // @[AxiLoadQueue.scala 131:41:@8711.4]
  assign _T_7682 = _T_7680 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8712.4]
  assign storesToCheck_0_2 = _T_2234 ? _T_7675 : _T_7682; // @[AxiLoadQueue.scala 130:10:@8713.4]
  assign _T_7688 = 4'h3 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8716.4]
  assign _T_7689 = _T_6172 & _T_7688; // @[AxiLoadQueue.scala 130:72:@8717.4]
  assign _T_7691 = offsetQ_0 < 4'h3; // @[AxiLoadQueue.scala 131:33:@8718.4]
  assign _T_7694 = _T_7691 & _T_6181; // @[AxiLoadQueue.scala 131:41:@8720.4]
  assign _T_7696 = _T_7694 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8721.4]
  assign storesToCheck_0_3 = _T_2234 ? _T_7689 : _T_7696; // @[AxiLoadQueue.scala 130:10:@8722.4]
  assign _T_7702 = 4'h4 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8725.4]
  assign _T_7703 = _T_6189 & _T_7702; // @[AxiLoadQueue.scala 130:72:@8726.4]
  assign _T_7705 = offsetQ_0 < 4'h4; // @[AxiLoadQueue.scala 131:33:@8727.4]
  assign _T_7708 = _T_7705 & _T_6198; // @[AxiLoadQueue.scala 131:41:@8729.4]
  assign _T_7710 = _T_7708 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8730.4]
  assign storesToCheck_0_4 = _T_2234 ? _T_7703 : _T_7710; // @[AxiLoadQueue.scala 130:10:@8731.4]
  assign _T_7716 = 4'h5 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8734.4]
  assign _T_7717 = _T_6206 & _T_7716; // @[AxiLoadQueue.scala 130:72:@8735.4]
  assign _T_7719 = offsetQ_0 < 4'h5; // @[AxiLoadQueue.scala 131:33:@8736.4]
  assign _T_7722 = _T_7719 & _T_6215; // @[AxiLoadQueue.scala 131:41:@8738.4]
  assign _T_7724 = _T_7722 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8739.4]
  assign storesToCheck_0_5 = _T_2234 ? _T_7717 : _T_7724; // @[AxiLoadQueue.scala 130:10:@8740.4]
  assign _T_7730 = 4'h6 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8743.4]
  assign _T_7731 = _T_6223 & _T_7730; // @[AxiLoadQueue.scala 130:72:@8744.4]
  assign _T_7733 = offsetQ_0 < 4'h6; // @[AxiLoadQueue.scala 131:33:@8745.4]
  assign _T_7736 = _T_7733 & _T_6232; // @[AxiLoadQueue.scala 131:41:@8747.4]
  assign _T_7738 = _T_7736 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8748.4]
  assign storesToCheck_0_6 = _T_2234 ? _T_7731 : _T_7738; // @[AxiLoadQueue.scala 130:10:@8749.4]
  assign _T_7744 = 4'h7 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8752.4]
  assign _T_7745 = _T_6240 & _T_7744; // @[AxiLoadQueue.scala 130:72:@8753.4]
  assign _T_7747 = offsetQ_0 < 4'h7; // @[AxiLoadQueue.scala 131:33:@8754.4]
  assign _T_7750 = _T_7747 & _T_6249; // @[AxiLoadQueue.scala 131:41:@8756.4]
  assign _T_7752 = _T_7750 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8757.4]
  assign storesToCheck_0_7 = _T_2234 ? _T_7745 : _T_7752; // @[AxiLoadQueue.scala 130:10:@8758.4]
  assign _T_7758 = 4'h8 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8761.4]
  assign _T_7759 = _T_6257 & _T_7758; // @[AxiLoadQueue.scala 130:72:@8762.4]
  assign _T_7761 = offsetQ_0 < 4'h8; // @[AxiLoadQueue.scala 131:33:@8763.4]
  assign _T_7764 = _T_7761 & _T_6266; // @[AxiLoadQueue.scala 131:41:@8765.4]
  assign _T_7766 = _T_7764 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8766.4]
  assign storesToCheck_0_8 = _T_2234 ? _T_7759 : _T_7766; // @[AxiLoadQueue.scala 130:10:@8767.4]
  assign _T_7772 = 4'h9 <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8770.4]
  assign _T_7773 = _T_6274 & _T_7772; // @[AxiLoadQueue.scala 130:72:@8771.4]
  assign _T_7775 = offsetQ_0 < 4'h9; // @[AxiLoadQueue.scala 131:33:@8772.4]
  assign _T_7778 = _T_7775 & _T_6283; // @[AxiLoadQueue.scala 131:41:@8774.4]
  assign _T_7780 = _T_7778 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8775.4]
  assign storesToCheck_0_9 = _T_2234 ? _T_7773 : _T_7780; // @[AxiLoadQueue.scala 130:10:@8776.4]
  assign _T_7786 = 4'ha <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8779.4]
  assign _T_7787 = _T_6291 & _T_7786; // @[AxiLoadQueue.scala 130:72:@8780.4]
  assign _T_7789 = offsetQ_0 < 4'ha; // @[AxiLoadQueue.scala 131:33:@8781.4]
  assign _T_7792 = _T_7789 & _T_6300; // @[AxiLoadQueue.scala 131:41:@8783.4]
  assign _T_7794 = _T_7792 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8784.4]
  assign storesToCheck_0_10 = _T_2234 ? _T_7787 : _T_7794; // @[AxiLoadQueue.scala 130:10:@8785.4]
  assign _T_7800 = 4'hb <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8788.4]
  assign _T_7801 = _T_6308 & _T_7800; // @[AxiLoadQueue.scala 130:72:@8789.4]
  assign _T_7803 = offsetQ_0 < 4'hb; // @[AxiLoadQueue.scala 131:33:@8790.4]
  assign _T_7806 = _T_7803 & _T_6317; // @[AxiLoadQueue.scala 131:41:@8792.4]
  assign _T_7808 = _T_7806 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8793.4]
  assign storesToCheck_0_11 = _T_2234 ? _T_7801 : _T_7808; // @[AxiLoadQueue.scala 130:10:@8794.4]
  assign _T_7814 = 4'hc <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8797.4]
  assign _T_7815 = _T_6325 & _T_7814; // @[AxiLoadQueue.scala 130:72:@8798.4]
  assign _T_7817 = offsetQ_0 < 4'hc; // @[AxiLoadQueue.scala 131:33:@8799.4]
  assign _T_7820 = _T_7817 & _T_6334; // @[AxiLoadQueue.scala 131:41:@8801.4]
  assign _T_7822 = _T_7820 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8802.4]
  assign storesToCheck_0_12 = _T_2234 ? _T_7815 : _T_7822; // @[AxiLoadQueue.scala 130:10:@8803.4]
  assign _T_7828 = 4'hd <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8806.4]
  assign _T_7829 = _T_6342 & _T_7828; // @[AxiLoadQueue.scala 130:72:@8807.4]
  assign _T_7831 = offsetQ_0 < 4'hd; // @[AxiLoadQueue.scala 131:33:@8808.4]
  assign _T_7834 = _T_7831 & _T_6351; // @[AxiLoadQueue.scala 131:41:@8810.4]
  assign _T_7836 = _T_7834 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8811.4]
  assign storesToCheck_0_13 = _T_2234 ? _T_7829 : _T_7836; // @[AxiLoadQueue.scala 130:10:@8812.4]
  assign _T_7842 = 4'he <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8815.4]
  assign _T_7843 = _T_6359 & _T_7842; // @[AxiLoadQueue.scala 130:72:@8816.4]
  assign _T_7845 = offsetQ_0 < 4'he; // @[AxiLoadQueue.scala 131:33:@8817.4]
  assign _T_7848 = _T_7845 & _T_6368; // @[AxiLoadQueue.scala 131:41:@8819.4]
  assign _T_7850 = _T_7848 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8820.4]
  assign storesToCheck_0_14 = _T_2234 ? _T_7843 : _T_7850; // @[AxiLoadQueue.scala 130:10:@8821.4]
  assign _T_7856 = 4'hf <= offsetQ_0; // @[AxiLoadQueue.scala 130:81:@8824.4]
  assign storesToCheck_0_15 = _T_2234 ? _T_7856 : 1'h1; // @[AxiLoadQueue.scala 130:10:@8830.4]
  assign storesToCheck_1_0 = _T_2264 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@8872.4]
  assign _T_7906 = 4'h1 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8875.4]
  assign _T_7907 = _T_6138 & _T_7906; // @[AxiLoadQueue.scala 130:72:@8876.4]
  assign _T_7909 = offsetQ_1 < 4'h1; // @[AxiLoadQueue.scala 131:33:@8877.4]
  assign _T_7912 = _T_7909 & _T_6147; // @[AxiLoadQueue.scala 131:41:@8879.4]
  assign _T_7914 = _T_7912 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8880.4]
  assign storesToCheck_1_1 = _T_2264 ? _T_7907 : _T_7914; // @[AxiLoadQueue.scala 130:10:@8881.4]
  assign _T_7920 = 4'h2 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8884.4]
  assign _T_7921 = _T_6155 & _T_7920; // @[AxiLoadQueue.scala 130:72:@8885.4]
  assign _T_7923 = offsetQ_1 < 4'h2; // @[AxiLoadQueue.scala 131:33:@8886.4]
  assign _T_7926 = _T_7923 & _T_6164; // @[AxiLoadQueue.scala 131:41:@8888.4]
  assign _T_7928 = _T_7926 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8889.4]
  assign storesToCheck_1_2 = _T_2264 ? _T_7921 : _T_7928; // @[AxiLoadQueue.scala 130:10:@8890.4]
  assign _T_7934 = 4'h3 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8893.4]
  assign _T_7935 = _T_6172 & _T_7934; // @[AxiLoadQueue.scala 130:72:@8894.4]
  assign _T_7937 = offsetQ_1 < 4'h3; // @[AxiLoadQueue.scala 131:33:@8895.4]
  assign _T_7940 = _T_7937 & _T_6181; // @[AxiLoadQueue.scala 131:41:@8897.4]
  assign _T_7942 = _T_7940 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8898.4]
  assign storesToCheck_1_3 = _T_2264 ? _T_7935 : _T_7942; // @[AxiLoadQueue.scala 130:10:@8899.4]
  assign _T_7948 = 4'h4 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8902.4]
  assign _T_7949 = _T_6189 & _T_7948; // @[AxiLoadQueue.scala 130:72:@8903.4]
  assign _T_7951 = offsetQ_1 < 4'h4; // @[AxiLoadQueue.scala 131:33:@8904.4]
  assign _T_7954 = _T_7951 & _T_6198; // @[AxiLoadQueue.scala 131:41:@8906.4]
  assign _T_7956 = _T_7954 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8907.4]
  assign storesToCheck_1_4 = _T_2264 ? _T_7949 : _T_7956; // @[AxiLoadQueue.scala 130:10:@8908.4]
  assign _T_7962 = 4'h5 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8911.4]
  assign _T_7963 = _T_6206 & _T_7962; // @[AxiLoadQueue.scala 130:72:@8912.4]
  assign _T_7965 = offsetQ_1 < 4'h5; // @[AxiLoadQueue.scala 131:33:@8913.4]
  assign _T_7968 = _T_7965 & _T_6215; // @[AxiLoadQueue.scala 131:41:@8915.4]
  assign _T_7970 = _T_7968 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8916.4]
  assign storesToCheck_1_5 = _T_2264 ? _T_7963 : _T_7970; // @[AxiLoadQueue.scala 130:10:@8917.4]
  assign _T_7976 = 4'h6 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8920.4]
  assign _T_7977 = _T_6223 & _T_7976; // @[AxiLoadQueue.scala 130:72:@8921.4]
  assign _T_7979 = offsetQ_1 < 4'h6; // @[AxiLoadQueue.scala 131:33:@8922.4]
  assign _T_7982 = _T_7979 & _T_6232; // @[AxiLoadQueue.scala 131:41:@8924.4]
  assign _T_7984 = _T_7982 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8925.4]
  assign storesToCheck_1_6 = _T_2264 ? _T_7977 : _T_7984; // @[AxiLoadQueue.scala 130:10:@8926.4]
  assign _T_7990 = 4'h7 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8929.4]
  assign _T_7991 = _T_6240 & _T_7990; // @[AxiLoadQueue.scala 130:72:@8930.4]
  assign _T_7993 = offsetQ_1 < 4'h7; // @[AxiLoadQueue.scala 131:33:@8931.4]
  assign _T_7996 = _T_7993 & _T_6249; // @[AxiLoadQueue.scala 131:41:@8933.4]
  assign _T_7998 = _T_7996 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8934.4]
  assign storesToCheck_1_7 = _T_2264 ? _T_7991 : _T_7998; // @[AxiLoadQueue.scala 130:10:@8935.4]
  assign _T_8004 = 4'h8 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8938.4]
  assign _T_8005 = _T_6257 & _T_8004; // @[AxiLoadQueue.scala 130:72:@8939.4]
  assign _T_8007 = offsetQ_1 < 4'h8; // @[AxiLoadQueue.scala 131:33:@8940.4]
  assign _T_8010 = _T_8007 & _T_6266; // @[AxiLoadQueue.scala 131:41:@8942.4]
  assign _T_8012 = _T_8010 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8943.4]
  assign storesToCheck_1_8 = _T_2264 ? _T_8005 : _T_8012; // @[AxiLoadQueue.scala 130:10:@8944.4]
  assign _T_8018 = 4'h9 <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8947.4]
  assign _T_8019 = _T_6274 & _T_8018; // @[AxiLoadQueue.scala 130:72:@8948.4]
  assign _T_8021 = offsetQ_1 < 4'h9; // @[AxiLoadQueue.scala 131:33:@8949.4]
  assign _T_8024 = _T_8021 & _T_6283; // @[AxiLoadQueue.scala 131:41:@8951.4]
  assign _T_8026 = _T_8024 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8952.4]
  assign storesToCheck_1_9 = _T_2264 ? _T_8019 : _T_8026; // @[AxiLoadQueue.scala 130:10:@8953.4]
  assign _T_8032 = 4'ha <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8956.4]
  assign _T_8033 = _T_6291 & _T_8032; // @[AxiLoadQueue.scala 130:72:@8957.4]
  assign _T_8035 = offsetQ_1 < 4'ha; // @[AxiLoadQueue.scala 131:33:@8958.4]
  assign _T_8038 = _T_8035 & _T_6300; // @[AxiLoadQueue.scala 131:41:@8960.4]
  assign _T_8040 = _T_8038 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8961.4]
  assign storesToCheck_1_10 = _T_2264 ? _T_8033 : _T_8040; // @[AxiLoadQueue.scala 130:10:@8962.4]
  assign _T_8046 = 4'hb <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8965.4]
  assign _T_8047 = _T_6308 & _T_8046; // @[AxiLoadQueue.scala 130:72:@8966.4]
  assign _T_8049 = offsetQ_1 < 4'hb; // @[AxiLoadQueue.scala 131:33:@8967.4]
  assign _T_8052 = _T_8049 & _T_6317; // @[AxiLoadQueue.scala 131:41:@8969.4]
  assign _T_8054 = _T_8052 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8970.4]
  assign storesToCheck_1_11 = _T_2264 ? _T_8047 : _T_8054; // @[AxiLoadQueue.scala 130:10:@8971.4]
  assign _T_8060 = 4'hc <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8974.4]
  assign _T_8061 = _T_6325 & _T_8060; // @[AxiLoadQueue.scala 130:72:@8975.4]
  assign _T_8063 = offsetQ_1 < 4'hc; // @[AxiLoadQueue.scala 131:33:@8976.4]
  assign _T_8066 = _T_8063 & _T_6334; // @[AxiLoadQueue.scala 131:41:@8978.4]
  assign _T_8068 = _T_8066 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8979.4]
  assign storesToCheck_1_12 = _T_2264 ? _T_8061 : _T_8068; // @[AxiLoadQueue.scala 130:10:@8980.4]
  assign _T_8074 = 4'hd <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8983.4]
  assign _T_8075 = _T_6342 & _T_8074; // @[AxiLoadQueue.scala 130:72:@8984.4]
  assign _T_8077 = offsetQ_1 < 4'hd; // @[AxiLoadQueue.scala 131:33:@8985.4]
  assign _T_8080 = _T_8077 & _T_6351; // @[AxiLoadQueue.scala 131:41:@8987.4]
  assign _T_8082 = _T_8080 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8988.4]
  assign storesToCheck_1_13 = _T_2264 ? _T_8075 : _T_8082; // @[AxiLoadQueue.scala 130:10:@8989.4]
  assign _T_8088 = 4'he <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@8992.4]
  assign _T_8089 = _T_6359 & _T_8088; // @[AxiLoadQueue.scala 130:72:@8993.4]
  assign _T_8091 = offsetQ_1 < 4'he; // @[AxiLoadQueue.scala 131:33:@8994.4]
  assign _T_8094 = _T_8091 & _T_6368; // @[AxiLoadQueue.scala 131:41:@8996.4]
  assign _T_8096 = _T_8094 == 1'h0; // @[AxiLoadQueue.scala 131:9:@8997.4]
  assign storesToCheck_1_14 = _T_2264 ? _T_8089 : _T_8096; // @[AxiLoadQueue.scala 130:10:@8998.4]
  assign _T_8102 = 4'hf <= offsetQ_1; // @[AxiLoadQueue.scala 130:81:@9001.4]
  assign storesToCheck_1_15 = _T_2264 ? _T_8102 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9007.4]
  assign storesToCheck_2_0 = _T_2294 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9049.4]
  assign _T_8152 = 4'h1 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9052.4]
  assign _T_8153 = _T_6138 & _T_8152; // @[AxiLoadQueue.scala 130:72:@9053.4]
  assign _T_8155 = offsetQ_2 < 4'h1; // @[AxiLoadQueue.scala 131:33:@9054.4]
  assign _T_8158 = _T_8155 & _T_6147; // @[AxiLoadQueue.scala 131:41:@9056.4]
  assign _T_8160 = _T_8158 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9057.4]
  assign storesToCheck_2_1 = _T_2294 ? _T_8153 : _T_8160; // @[AxiLoadQueue.scala 130:10:@9058.4]
  assign _T_8166 = 4'h2 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9061.4]
  assign _T_8167 = _T_6155 & _T_8166; // @[AxiLoadQueue.scala 130:72:@9062.4]
  assign _T_8169 = offsetQ_2 < 4'h2; // @[AxiLoadQueue.scala 131:33:@9063.4]
  assign _T_8172 = _T_8169 & _T_6164; // @[AxiLoadQueue.scala 131:41:@9065.4]
  assign _T_8174 = _T_8172 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9066.4]
  assign storesToCheck_2_2 = _T_2294 ? _T_8167 : _T_8174; // @[AxiLoadQueue.scala 130:10:@9067.4]
  assign _T_8180 = 4'h3 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9070.4]
  assign _T_8181 = _T_6172 & _T_8180; // @[AxiLoadQueue.scala 130:72:@9071.4]
  assign _T_8183 = offsetQ_2 < 4'h3; // @[AxiLoadQueue.scala 131:33:@9072.4]
  assign _T_8186 = _T_8183 & _T_6181; // @[AxiLoadQueue.scala 131:41:@9074.4]
  assign _T_8188 = _T_8186 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9075.4]
  assign storesToCheck_2_3 = _T_2294 ? _T_8181 : _T_8188; // @[AxiLoadQueue.scala 130:10:@9076.4]
  assign _T_8194 = 4'h4 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9079.4]
  assign _T_8195 = _T_6189 & _T_8194; // @[AxiLoadQueue.scala 130:72:@9080.4]
  assign _T_8197 = offsetQ_2 < 4'h4; // @[AxiLoadQueue.scala 131:33:@9081.4]
  assign _T_8200 = _T_8197 & _T_6198; // @[AxiLoadQueue.scala 131:41:@9083.4]
  assign _T_8202 = _T_8200 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9084.4]
  assign storesToCheck_2_4 = _T_2294 ? _T_8195 : _T_8202; // @[AxiLoadQueue.scala 130:10:@9085.4]
  assign _T_8208 = 4'h5 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9088.4]
  assign _T_8209 = _T_6206 & _T_8208; // @[AxiLoadQueue.scala 130:72:@9089.4]
  assign _T_8211 = offsetQ_2 < 4'h5; // @[AxiLoadQueue.scala 131:33:@9090.4]
  assign _T_8214 = _T_8211 & _T_6215; // @[AxiLoadQueue.scala 131:41:@9092.4]
  assign _T_8216 = _T_8214 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9093.4]
  assign storesToCheck_2_5 = _T_2294 ? _T_8209 : _T_8216; // @[AxiLoadQueue.scala 130:10:@9094.4]
  assign _T_8222 = 4'h6 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9097.4]
  assign _T_8223 = _T_6223 & _T_8222; // @[AxiLoadQueue.scala 130:72:@9098.4]
  assign _T_8225 = offsetQ_2 < 4'h6; // @[AxiLoadQueue.scala 131:33:@9099.4]
  assign _T_8228 = _T_8225 & _T_6232; // @[AxiLoadQueue.scala 131:41:@9101.4]
  assign _T_8230 = _T_8228 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9102.4]
  assign storesToCheck_2_6 = _T_2294 ? _T_8223 : _T_8230; // @[AxiLoadQueue.scala 130:10:@9103.4]
  assign _T_8236 = 4'h7 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9106.4]
  assign _T_8237 = _T_6240 & _T_8236; // @[AxiLoadQueue.scala 130:72:@9107.4]
  assign _T_8239 = offsetQ_2 < 4'h7; // @[AxiLoadQueue.scala 131:33:@9108.4]
  assign _T_8242 = _T_8239 & _T_6249; // @[AxiLoadQueue.scala 131:41:@9110.4]
  assign _T_8244 = _T_8242 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9111.4]
  assign storesToCheck_2_7 = _T_2294 ? _T_8237 : _T_8244; // @[AxiLoadQueue.scala 130:10:@9112.4]
  assign _T_8250 = 4'h8 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9115.4]
  assign _T_8251 = _T_6257 & _T_8250; // @[AxiLoadQueue.scala 130:72:@9116.4]
  assign _T_8253 = offsetQ_2 < 4'h8; // @[AxiLoadQueue.scala 131:33:@9117.4]
  assign _T_8256 = _T_8253 & _T_6266; // @[AxiLoadQueue.scala 131:41:@9119.4]
  assign _T_8258 = _T_8256 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9120.4]
  assign storesToCheck_2_8 = _T_2294 ? _T_8251 : _T_8258; // @[AxiLoadQueue.scala 130:10:@9121.4]
  assign _T_8264 = 4'h9 <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9124.4]
  assign _T_8265 = _T_6274 & _T_8264; // @[AxiLoadQueue.scala 130:72:@9125.4]
  assign _T_8267 = offsetQ_2 < 4'h9; // @[AxiLoadQueue.scala 131:33:@9126.4]
  assign _T_8270 = _T_8267 & _T_6283; // @[AxiLoadQueue.scala 131:41:@9128.4]
  assign _T_8272 = _T_8270 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9129.4]
  assign storesToCheck_2_9 = _T_2294 ? _T_8265 : _T_8272; // @[AxiLoadQueue.scala 130:10:@9130.4]
  assign _T_8278 = 4'ha <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9133.4]
  assign _T_8279 = _T_6291 & _T_8278; // @[AxiLoadQueue.scala 130:72:@9134.4]
  assign _T_8281 = offsetQ_2 < 4'ha; // @[AxiLoadQueue.scala 131:33:@9135.4]
  assign _T_8284 = _T_8281 & _T_6300; // @[AxiLoadQueue.scala 131:41:@9137.4]
  assign _T_8286 = _T_8284 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9138.4]
  assign storesToCheck_2_10 = _T_2294 ? _T_8279 : _T_8286; // @[AxiLoadQueue.scala 130:10:@9139.4]
  assign _T_8292 = 4'hb <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9142.4]
  assign _T_8293 = _T_6308 & _T_8292; // @[AxiLoadQueue.scala 130:72:@9143.4]
  assign _T_8295 = offsetQ_2 < 4'hb; // @[AxiLoadQueue.scala 131:33:@9144.4]
  assign _T_8298 = _T_8295 & _T_6317; // @[AxiLoadQueue.scala 131:41:@9146.4]
  assign _T_8300 = _T_8298 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9147.4]
  assign storesToCheck_2_11 = _T_2294 ? _T_8293 : _T_8300; // @[AxiLoadQueue.scala 130:10:@9148.4]
  assign _T_8306 = 4'hc <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9151.4]
  assign _T_8307 = _T_6325 & _T_8306; // @[AxiLoadQueue.scala 130:72:@9152.4]
  assign _T_8309 = offsetQ_2 < 4'hc; // @[AxiLoadQueue.scala 131:33:@9153.4]
  assign _T_8312 = _T_8309 & _T_6334; // @[AxiLoadQueue.scala 131:41:@9155.4]
  assign _T_8314 = _T_8312 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9156.4]
  assign storesToCheck_2_12 = _T_2294 ? _T_8307 : _T_8314; // @[AxiLoadQueue.scala 130:10:@9157.4]
  assign _T_8320 = 4'hd <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9160.4]
  assign _T_8321 = _T_6342 & _T_8320; // @[AxiLoadQueue.scala 130:72:@9161.4]
  assign _T_8323 = offsetQ_2 < 4'hd; // @[AxiLoadQueue.scala 131:33:@9162.4]
  assign _T_8326 = _T_8323 & _T_6351; // @[AxiLoadQueue.scala 131:41:@9164.4]
  assign _T_8328 = _T_8326 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9165.4]
  assign storesToCheck_2_13 = _T_2294 ? _T_8321 : _T_8328; // @[AxiLoadQueue.scala 130:10:@9166.4]
  assign _T_8334 = 4'he <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9169.4]
  assign _T_8335 = _T_6359 & _T_8334; // @[AxiLoadQueue.scala 130:72:@9170.4]
  assign _T_8337 = offsetQ_2 < 4'he; // @[AxiLoadQueue.scala 131:33:@9171.4]
  assign _T_8340 = _T_8337 & _T_6368; // @[AxiLoadQueue.scala 131:41:@9173.4]
  assign _T_8342 = _T_8340 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9174.4]
  assign storesToCheck_2_14 = _T_2294 ? _T_8335 : _T_8342; // @[AxiLoadQueue.scala 130:10:@9175.4]
  assign _T_8348 = 4'hf <= offsetQ_2; // @[AxiLoadQueue.scala 130:81:@9178.4]
  assign storesToCheck_2_15 = _T_2294 ? _T_8348 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9184.4]
  assign storesToCheck_3_0 = _T_2324 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9226.4]
  assign _T_8398 = 4'h1 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9229.4]
  assign _T_8399 = _T_6138 & _T_8398; // @[AxiLoadQueue.scala 130:72:@9230.4]
  assign _T_8401 = offsetQ_3 < 4'h1; // @[AxiLoadQueue.scala 131:33:@9231.4]
  assign _T_8404 = _T_8401 & _T_6147; // @[AxiLoadQueue.scala 131:41:@9233.4]
  assign _T_8406 = _T_8404 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9234.4]
  assign storesToCheck_3_1 = _T_2324 ? _T_8399 : _T_8406; // @[AxiLoadQueue.scala 130:10:@9235.4]
  assign _T_8412 = 4'h2 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9238.4]
  assign _T_8413 = _T_6155 & _T_8412; // @[AxiLoadQueue.scala 130:72:@9239.4]
  assign _T_8415 = offsetQ_3 < 4'h2; // @[AxiLoadQueue.scala 131:33:@9240.4]
  assign _T_8418 = _T_8415 & _T_6164; // @[AxiLoadQueue.scala 131:41:@9242.4]
  assign _T_8420 = _T_8418 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9243.4]
  assign storesToCheck_3_2 = _T_2324 ? _T_8413 : _T_8420; // @[AxiLoadQueue.scala 130:10:@9244.4]
  assign _T_8426 = 4'h3 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9247.4]
  assign _T_8427 = _T_6172 & _T_8426; // @[AxiLoadQueue.scala 130:72:@9248.4]
  assign _T_8429 = offsetQ_3 < 4'h3; // @[AxiLoadQueue.scala 131:33:@9249.4]
  assign _T_8432 = _T_8429 & _T_6181; // @[AxiLoadQueue.scala 131:41:@9251.4]
  assign _T_8434 = _T_8432 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9252.4]
  assign storesToCheck_3_3 = _T_2324 ? _T_8427 : _T_8434; // @[AxiLoadQueue.scala 130:10:@9253.4]
  assign _T_8440 = 4'h4 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9256.4]
  assign _T_8441 = _T_6189 & _T_8440; // @[AxiLoadQueue.scala 130:72:@9257.4]
  assign _T_8443 = offsetQ_3 < 4'h4; // @[AxiLoadQueue.scala 131:33:@9258.4]
  assign _T_8446 = _T_8443 & _T_6198; // @[AxiLoadQueue.scala 131:41:@9260.4]
  assign _T_8448 = _T_8446 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9261.4]
  assign storesToCheck_3_4 = _T_2324 ? _T_8441 : _T_8448; // @[AxiLoadQueue.scala 130:10:@9262.4]
  assign _T_8454 = 4'h5 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9265.4]
  assign _T_8455 = _T_6206 & _T_8454; // @[AxiLoadQueue.scala 130:72:@9266.4]
  assign _T_8457 = offsetQ_3 < 4'h5; // @[AxiLoadQueue.scala 131:33:@9267.4]
  assign _T_8460 = _T_8457 & _T_6215; // @[AxiLoadQueue.scala 131:41:@9269.4]
  assign _T_8462 = _T_8460 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9270.4]
  assign storesToCheck_3_5 = _T_2324 ? _T_8455 : _T_8462; // @[AxiLoadQueue.scala 130:10:@9271.4]
  assign _T_8468 = 4'h6 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9274.4]
  assign _T_8469 = _T_6223 & _T_8468; // @[AxiLoadQueue.scala 130:72:@9275.4]
  assign _T_8471 = offsetQ_3 < 4'h6; // @[AxiLoadQueue.scala 131:33:@9276.4]
  assign _T_8474 = _T_8471 & _T_6232; // @[AxiLoadQueue.scala 131:41:@9278.4]
  assign _T_8476 = _T_8474 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9279.4]
  assign storesToCheck_3_6 = _T_2324 ? _T_8469 : _T_8476; // @[AxiLoadQueue.scala 130:10:@9280.4]
  assign _T_8482 = 4'h7 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9283.4]
  assign _T_8483 = _T_6240 & _T_8482; // @[AxiLoadQueue.scala 130:72:@9284.4]
  assign _T_8485 = offsetQ_3 < 4'h7; // @[AxiLoadQueue.scala 131:33:@9285.4]
  assign _T_8488 = _T_8485 & _T_6249; // @[AxiLoadQueue.scala 131:41:@9287.4]
  assign _T_8490 = _T_8488 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9288.4]
  assign storesToCheck_3_7 = _T_2324 ? _T_8483 : _T_8490; // @[AxiLoadQueue.scala 130:10:@9289.4]
  assign _T_8496 = 4'h8 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9292.4]
  assign _T_8497 = _T_6257 & _T_8496; // @[AxiLoadQueue.scala 130:72:@9293.4]
  assign _T_8499 = offsetQ_3 < 4'h8; // @[AxiLoadQueue.scala 131:33:@9294.4]
  assign _T_8502 = _T_8499 & _T_6266; // @[AxiLoadQueue.scala 131:41:@9296.4]
  assign _T_8504 = _T_8502 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9297.4]
  assign storesToCheck_3_8 = _T_2324 ? _T_8497 : _T_8504; // @[AxiLoadQueue.scala 130:10:@9298.4]
  assign _T_8510 = 4'h9 <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9301.4]
  assign _T_8511 = _T_6274 & _T_8510; // @[AxiLoadQueue.scala 130:72:@9302.4]
  assign _T_8513 = offsetQ_3 < 4'h9; // @[AxiLoadQueue.scala 131:33:@9303.4]
  assign _T_8516 = _T_8513 & _T_6283; // @[AxiLoadQueue.scala 131:41:@9305.4]
  assign _T_8518 = _T_8516 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9306.4]
  assign storesToCheck_3_9 = _T_2324 ? _T_8511 : _T_8518; // @[AxiLoadQueue.scala 130:10:@9307.4]
  assign _T_8524 = 4'ha <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9310.4]
  assign _T_8525 = _T_6291 & _T_8524; // @[AxiLoadQueue.scala 130:72:@9311.4]
  assign _T_8527 = offsetQ_3 < 4'ha; // @[AxiLoadQueue.scala 131:33:@9312.4]
  assign _T_8530 = _T_8527 & _T_6300; // @[AxiLoadQueue.scala 131:41:@9314.4]
  assign _T_8532 = _T_8530 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9315.4]
  assign storesToCheck_3_10 = _T_2324 ? _T_8525 : _T_8532; // @[AxiLoadQueue.scala 130:10:@9316.4]
  assign _T_8538 = 4'hb <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9319.4]
  assign _T_8539 = _T_6308 & _T_8538; // @[AxiLoadQueue.scala 130:72:@9320.4]
  assign _T_8541 = offsetQ_3 < 4'hb; // @[AxiLoadQueue.scala 131:33:@9321.4]
  assign _T_8544 = _T_8541 & _T_6317; // @[AxiLoadQueue.scala 131:41:@9323.4]
  assign _T_8546 = _T_8544 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9324.4]
  assign storesToCheck_3_11 = _T_2324 ? _T_8539 : _T_8546; // @[AxiLoadQueue.scala 130:10:@9325.4]
  assign _T_8552 = 4'hc <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9328.4]
  assign _T_8553 = _T_6325 & _T_8552; // @[AxiLoadQueue.scala 130:72:@9329.4]
  assign _T_8555 = offsetQ_3 < 4'hc; // @[AxiLoadQueue.scala 131:33:@9330.4]
  assign _T_8558 = _T_8555 & _T_6334; // @[AxiLoadQueue.scala 131:41:@9332.4]
  assign _T_8560 = _T_8558 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9333.4]
  assign storesToCheck_3_12 = _T_2324 ? _T_8553 : _T_8560; // @[AxiLoadQueue.scala 130:10:@9334.4]
  assign _T_8566 = 4'hd <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9337.4]
  assign _T_8567 = _T_6342 & _T_8566; // @[AxiLoadQueue.scala 130:72:@9338.4]
  assign _T_8569 = offsetQ_3 < 4'hd; // @[AxiLoadQueue.scala 131:33:@9339.4]
  assign _T_8572 = _T_8569 & _T_6351; // @[AxiLoadQueue.scala 131:41:@9341.4]
  assign _T_8574 = _T_8572 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9342.4]
  assign storesToCheck_3_13 = _T_2324 ? _T_8567 : _T_8574; // @[AxiLoadQueue.scala 130:10:@9343.4]
  assign _T_8580 = 4'he <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9346.4]
  assign _T_8581 = _T_6359 & _T_8580; // @[AxiLoadQueue.scala 130:72:@9347.4]
  assign _T_8583 = offsetQ_3 < 4'he; // @[AxiLoadQueue.scala 131:33:@9348.4]
  assign _T_8586 = _T_8583 & _T_6368; // @[AxiLoadQueue.scala 131:41:@9350.4]
  assign _T_8588 = _T_8586 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9351.4]
  assign storesToCheck_3_14 = _T_2324 ? _T_8581 : _T_8588; // @[AxiLoadQueue.scala 130:10:@9352.4]
  assign _T_8594 = 4'hf <= offsetQ_3; // @[AxiLoadQueue.scala 130:81:@9355.4]
  assign storesToCheck_3_15 = _T_2324 ? _T_8594 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9361.4]
  assign storesToCheck_4_0 = _T_2354 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9403.4]
  assign _T_8644 = 4'h1 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9406.4]
  assign _T_8645 = _T_6138 & _T_8644; // @[AxiLoadQueue.scala 130:72:@9407.4]
  assign _T_8647 = offsetQ_4 < 4'h1; // @[AxiLoadQueue.scala 131:33:@9408.4]
  assign _T_8650 = _T_8647 & _T_6147; // @[AxiLoadQueue.scala 131:41:@9410.4]
  assign _T_8652 = _T_8650 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9411.4]
  assign storesToCheck_4_1 = _T_2354 ? _T_8645 : _T_8652; // @[AxiLoadQueue.scala 130:10:@9412.4]
  assign _T_8658 = 4'h2 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9415.4]
  assign _T_8659 = _T_6155 & _T_8658; // @[AxiLoadQueue.scala 130:72:@9416.4]
  assign _T_8661 = offsetQ_4 < 4'h2; // @[AxiLoadQueue.scala 131:33:@9417.4]
  assign _T_8664 = _T_8661 & _T_6164; // @[AxiLoadQueue.scala 131:41:@9419.4]
  assign _T_8666 = _T_8664 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9420.4]
  assign storesToCheck_4_2 = _T_2354 ? _T_8659 : _T_8666; // @[AxiLoadQueue.scala 130:10:@9421.4]
  assign _T_8672 = 4'h3 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9424.4]
  assign _T_8673 = _T_6172 & _T_8672; // @[AxiLoadQueue.scala 130:72:@9425.4]
  assign _T_8675 = offsetQ_4 < 4'h3; // @[AxiLoadQueue.scala 131:33:@9426.4]
  assign _T_8678 = _T_8675 & _T_6181; // @[AxiLoadQueue.scala 131:41:@9428.4]
  assign _T_8680 = _T_8678 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9429.4]
  assign storesToCheck_4_3 = _T_2354 ? _T_8673 : _T_8680; // @[AxiLoadQueue.scala 130:10:@9430.4]
  assign _T_8686 = 4'h4 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9433.4]
  assign _T_8687 = _T_6189 & _T_8686; // @[AxiLoadQueue.scala 130:72:@9434.4]
  assign _T_8689 = offsetQ_4 < 4'h4; // @[AxiLoadQueue.scala 131:33:@9435.4]
  assign _T_8692 = _T_8689 & _T_6198; // @[AxiLoadQueue.scala 131:41:@9437.4]
  assign _T_8694 = _T_8692 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9438.4]
  assign storesToCheck_4_4 = _T_2354 ? _T_8687 : _T_8694; // @[AxiLoadQueue.scala 130:10:@9439.4]
  assign _T_8700 = 4'h5 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9442.4]
  assign _T_8701 = _T_6206 & _T_8700; // @[AxiLoadQueue.scala 130:72:@9443.4]
  assign _T_8703 = offsetQ_4 < 4'h5; // @[AxiLoadQueue.scala 131:33:@9444.4]
  assign _T_8706 = _T_8703 & _T_6215; // @[AxiLoadQueue.scala 131:41:@9446.4]
  assign _T_8708 = _T_8706 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9447.4]
  assign storesToCheck_4_5 = _T_2354 ? _T_8701 : _T_8708; // @[AxiLoadQueue.scala 130:10:@9448.4]
  assign _T_8714 = 4'h6 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9451.4]
  assign _T_8715 = _T_6223 & _T_8714; // @[AxiLoadQueue.scala 130:72:@9452.4]
  assign _T_8717 = offsetQ_4 < 4'h6; // @[AxiLoadQueue.scala 131:33:@9453.4]
  assign _T_8720 = _T_8717 & _T_6232; // @[AxiLoadQueue.scala 131:41:@9455.4]
  assign _T_8722 = _T_8720 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9456.4]
  assign storesToCheck_4_6 = _T_2354 ? _T_8715 : _T_8722; // @[AxiLoadQueue.scala 130:10:@9457.4]
  assign _T_8728 = 4'h7 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9460.4]
  assign _T_8729 = _T_6240 & _T_8728; // @[AxiLoadQueue.scala 130:72:@9461.4]
  assign _T_8731 = offsetQ_4 < 4'h7; // @[AxiLoadQueue.scala 131:33:@9462.4]
  assign _T_8734 = _T_8731 & _T_6249; // @[AxiLoadQueue.scala 131:41:@9464.4]
  assign _T_8736 = _T_8734 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9465.4]
  assign storesToCheck_4_7 = _T_2354 ? _T_8729 : _T_8736; // @[AxiLoadQueue.scala 130:10:@9466.4]
  assign _T_8742 = 4'h8 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9469.4]
  assign _T_8743 = _T_6257 & _T_8742; // @[AxiLoadQueue.scala 130:72:@9470.4]
  assign _T_8745 = offsetQ_4 < 4'h8; // @[AxiLoadQueue.scala 131:33:@9471.4]
  assign _T_8748 = _T_8745 & _T_6266; // @[AxiLoadQueue.scala 131:41:@9473.4]
  assign _T_8750 = _T_8748 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9474.4]
  assign storesToCheck_4_8 = _T_2354 ? _T_8743 : _T_8750; // @[AxiLoadQueue.scala 130:10:@9475.4]
  assign _T_8756 = 4'h9 <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9478.4]
  assign _T_8757 = _T_6274 & _T_8756; // @[AxiLoadQueue.scala 130:72:@9479.4]
  assign _T_8759 = offsetQ_4 < 4'h9; // @[AxiLoadQueue.scala 131:33:@9480.4]
  assign _T_8762 = _T_8759 & _T_6283; // @[AxiLoadQueue.scala 131:41:@9482.4]
  assign _T_8764 = _T_8762 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9483.4]
  assign storesToCheck_4_9 = _T_2354 ? _T_8757 : _T_8764; // @[AxiLoadQueue.scala 130:10:@9484.4]
  assign _T_8770 = 4'ha <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9487.4]
  assign _T_8771 = _T_6291 & _T_8770; // @[AxiLoadQueue.scala 130:72:@9488.4]
  assign _T_8773 = offsetQ_4 < 4'ha; // @[AxiLoadQueue.scala 131:33:@9489.4]
  assign _T_8776 = _T_8773 & _T_6300; // @[AxiLoadQueue.scala 131:41:@9491.4]
  assign _T_8778 = _T_8776 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9492.4]
  assign storesToCheck_4_10 = _T_2354 ? _T_8771 : _T_8778; // @[AxiLoadQueue.scala 130:10:@9493.4]
  assign _T_8784 = 4'hb <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9496.4]
  assign _T_8785 = _T_6308 & _T_8784; // @[AxiLoadQueue.scala 130:72:@9497.4]
  assign _T_8787 = offsetQ_4 < 4'hb; // @[AxiLoadQueue.scala 131:33:@9498.4]
  assign _T_8790 = _T_8787 & _T_6317; // @[AxiLoadQueue.scala 131:41:@9500.4]
  assign _T_8792 = _T_8790 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9501.4]
  assign storesToCheck_4_11 = _T_2354 ? _T_8785 : _T_8792; // @[AxiLoadQueue.scala 130:10:@9502.4]
  assign _T_8798 = 4'hc <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9505.4]
  assign _T_8799 = _T_6325 & _T_8798; // @[AxiLoadQueue.scala 130:72:@9506.4]
  assign _T_8801 = offsetQ_4 < 4'hc; // @[AxiLoadQueue.scala 131:33:@9507.4]
  assign _T_8804 = _T_8801 & _T_6334; // @[AxiLoadQueue.scala 131:41:@9509.4]
  assign _T_8806 = _T_8804 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9510.4]
  assign storesToCheck_4_12 = _T_2354 ? _T_8799 : _T_8806; // @[AxiLoadQueue.scala 130:10:@9511.4]
  assign _T_8812 = 4'hd <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9514.4]
  assign _T_8813 = _T_6342 & _T_8812; // @[AxiLoadQueue.scala 130:72:@9515.4]
  assign _T_8815 = offsetQ_4 < 4'hd; // @[AxiLoadQueue.scala 131:33:@9516.4]
  assign _T_8818 = _T_8815 & _T_6351; // @[AxiLoadQueue.scala 131:41:@9518.4]
  assign _T_8820 = _T_8818 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9519.4]
  assign storesToCheck_4_13 = _T_2354 ? _T_8813 : _T_8820; // @[AxiLoadQueue.scala 130:10:@9520.4]
  assign _T_8826 = 4'he <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9523.4]
  assign _T_8827 = _T_6359 & _T_8826; // @[AxiLoadQueue.scala 130:72:@9524.4]
  assign _T_8829 = offsetQ_4 < 4'he; // @[AxiLoadQueue.scala 131:33:@9525.4]
  assign _T_8832 = _T_8829 & _T_6368; // @[AxiLoadQueue.scala 131:41:@9527.4]
  assign _T_8834 = _T_8832 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9528.4]
  assign storesToCheck_4_14 = _T_2354 ? _T_8827 : _T_8834; // @[AxiLoadQueue.scala 130:10:@9529.4]
  assign _T_8840 = 4'hf <= offsetQ_4; // @[AxiLoadQueue.scala 130:81:@9532.4]
  assign storesToCheck_4_15 = _T_2354 ? _T_8840 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9538.4]
  assign storesToCheck_5_0 = _T_2384 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9580.4]
  assign _T_8890 = 4'h1 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9583.4]
  assign _T_8891 = _T_6138 & _T_8890; // @[AxiLoadQueue.scala 130:72:@9584.4]
  assign _T_8893 = offsetQ_5 < 4'h1; // @[AxiLoadQueue.scala 131:33:@9585.4]
  assign _T_8896 = _T_8893 & _T_6147; // @[AxiLoadQueue.scala 131:41:@9587.4]
  assign _T_8898 = _T_8896 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9588.4]
  assign storesToCheck_5_1 = _T_2384 ? _T_8891 : _T_8898; // @[AxiLoadQueue.scala 130:10:@9589.4]
  assign _T_8904 = 4'h2 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9592.4]
  assign _T_8905 = _T_6155 & _T_8904; // @[AxiLoadQueue.scala 130:72:@9593.4]
  assign _T_8907 = offsetQ_5 < 4'h2; // @[AxiLoadQueue.scala 131:33:@9594.4]
  assign _T_8910 = _T_8907 & _T_6164; // @[AxiLoadQueue.scala 131:41:@9596.4]
  assign _T_8912 = _T_8910 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9597.4]
  assign storesToCheck_5_2 = _T_2384 ? _T_8905 : _T_8912; // @[AxiLoadQueue.scala 130:10:@9598.4]
  assign _T_8918 = 4'h3 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9601.4]
  assign _T_8919 = _T_6172 & _T_8918; // @[AxiLoadQueue.scala 130:72:@9602.4]
  assign _T_8921 = offsetQ_5 < 4'h3; // @[AxiLoadQueue.scala 131:33:@9603.4]
  assign _T_8924 = _T_8921 & _T_6181; // @[AxiLoadQueue.scala 131:41:@9605.4]
  assign _T_8926 = _T_8924 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9606.4]
  assign storesToCheck_5_3 = _T_2384 ? _T_8919 : _T_8926; // @[AxiLoadQueue.scala 130:10:@9607.4]
  assign _T_8932 = 4'h4 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9610.4]
  assign _T_8933 = _T_6189 & _T_8932; // @[AxiLoadQueue.scala 130:72:@9611.4]
  assign _T_8935 = offsetQ_5 < 4'h4; // @[AxiLoadQueue.scala 131:33:@9612.4]
  assign _T_8938 = _T_8935 & _T_6198; // @[AxiLoadQueue.scala 131:41:@9614.4]
  assign _T_8940 = _T_8938 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9615.4]
  assign storesToCheck_5_4 = _T_2384 ? _T_8933 : _T_8940; // @[AxiLoadQueue.scala 130:10:@9616.4]
  assign _T_8946 = 4'h5 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9619.4]
  assign _T_8947 = _T_6206 & _T_8946; // @[AxiLoadQueue.scala 130:72:@9620.4]
  assign _T_8949 = offsetQ_5 < 4'h5; // @[AxiLoadQueue.scala 131:33:@9621.4]
  assign _T_8952 = _T_8949 & _T_6215; // @[AxiLoadQueue.scala 131:41:@9623.4]
  assign _T_8954 = _T_8952 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9624.4]
  assign storesToCheck_5_5 = _T_2384 ? _T_8947 : _T_8954; // @[AxiLoadQueue.scala 130:10:@9625.4]
  assign _T_8960 = 4'h6 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9628.4]
  assign _T_8961 = _T_6223 & _T_8960; // @[AxiLoadQueue.scala 130:72:@9629.4]
  assign _T_8963 = offsetQ_5 < 4'h6; // @[AxiLoadQueue.scala 131:33:@9630.4]
  assign _T_8966 = _T_8963 & _T_6232; // @[AxiLoadQueue.scala 131:41:@9632.4]
  assign _T_8968 = _T_8966 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9633.4]
  assign storesToCheck_5_6 = _T_2384 ? _T_8961 : _T_8968; // @[AxiLoadQueue.scala 130:10:@9634.4]
  assign _T_8974 = 4'h7 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9637.4]
  assign _T_8975 = _T_6240 & _T_8974; // @[AxiLoadQueue.scala 130:72:@9638.4]
  assign _T_8977 = offsetQ_5 < 4'h7; // @[AxiLoadQueue.scala 131:33:@9639.4]
  assign _T_8980 = _T_8977 & _T_6249; // @[AxiLoadQueue.scala 131:41:@9641.4]
  assign _T_8982 = _T_8980 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9642.4]
  assign storesToCheck_5_7 = _T_2384 ? _T_8975 : _T_8982; // @[AxiLoadQueue.scala 130:10:@9643.4]
  assign _T_8988 = 4'h8 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9646.4]
  assign _T_8989 = _T_6257 & _T_8988; // @[AxiLoadQueue.scala 130:72:@9647.4]
  assign _T_8991 = offsetQ_5 < 4'h8; // @[AxiLoadQueue.scala 131:33:@9648.4]
  assign _T_8994 = _T_8991 & _T_6266; // @[AxiLoadQueue.scala 131:41:@9650.4]
  assign _T_8996 = _T_8994 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9651.4]
  assign storesToCheck_5_8 = _T_2384 ? _T_8989 : _T_8996; // @[AxiLoadQueue.scala 130:10:@9652.4]
  assign _T_9002 = 4'h9 <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9655.4]
  assign _T_9003 = _T_6274 & _T_9002; // @[AxiLoadQueue.scala 130:72:@9656.4]
  assign _T_9005 = offsetQ_5 < 4'h9; // @[AxiLoadQueue.scala 131:33:@9657.4]
  assign _T_9008 = _T_9005 & _T_6283; // @[AxiLoadQueue.scala 131:41:@9659.4]
  assign _T_9010 = _T_9008 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9660.4]
  assign storesToCheck_5_9 = _T_2384 ? _T_9003 : _T_9010; // @[AxiLoadQueue.scala 130:10:@9661.4]
  assign _T_9016 = 4'ha <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9664.4]
  assign _T_9017 = _T_6291 & _T_9016; // @[AxiLoadQueue.scala 130:72:@9665.4]
  assign _T_9019 = offsetQ_5 < 4'ha; // @[AxiLoadQueue.scala 131:33:@9666.4]
  assign _T_9022 = _T_9019 & _T_6300; // @[AxiLoadQueue.scala 131:41:@9668.4]
  assign _T_9024 = _T_9022 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9669.4]
  assign storesToCheck_5_10 = _T_2384 ? _T_9017 : _T_9024; // @[AxiLoadQueue.scala 130:10:@9670.4]
  assign _T_9030 = 4'hb <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9673.4]
  assign _T_9031 = _T_6308 & _T_9030; // @[AxiLoadQueue.scala 130:72:@9674.4]
  assign _T_9033 = offsetQ_5 < 4'hb; // @[AxiLoadQueue.scala 131:33:@9675.4]
  assign _T_9036 = _T_9033 & _T_6317; // @[AxiLoadQueue.scala 131:41:@9677.4]
  assign _T_9038 = _T_9036 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9678.4]
  assign storesToCheck_5_11 = _T_2384 ? _T_9031 : _T_9038; // @[AxiLoadQueue.scala 130:10:@9679.4]
  assign _T_9044 = 4'hc <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9682.4]
  assign _T_9045 = _T_6325 & _T_9044; // @[AxiLoadQueue.scala 130:72:@9683.4]
  assign _T_9047 = offsetQ_5 < 4'hc; // @[AxiLoadQueue.scala 131:33:@9684.4]
  assign _T_9050 = _T_9047 & _T_6334; // @[AxiLoadQueue.scala 131:41:@9686.4]
  assign _T_9052 = _T_9050 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9687.4]
  assign storesToCheck_5_12 = _T_2384 ? _T_9045 : _T_9052; // @[AxiLoadQueue.scala 130:10:@9688.4]
  assign _T_9058 = 4'hd <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9691.4]
  assign _T_9059 = _T_6342 & _T_9058; // @[AxiLoadQueue.scala 130:72:@9692.4]
  assign _T_9061 = offsetQ_5 < 4'hd; // @[AxiLoadQueue.scala 131:33:@9693.4]
  assign _T_9064 = _T_9061 & _T_6351; // @[AxiLoadQueue.scala 131:41:@9695.4]
  assign _T_9066 = _T_9064 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9696.4]
  assign storesToCheck_5_13 = _T_2384 ? _T_9059 : _T_9066; // @[AxiLoadQueue.scala 130:10:@9697.4]
  assign _T_9072 = 4'he <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9700.4]
  assign _T_9073 = _T_6359 & _T_9072; // @[AxiLoadQueue.scala 130:72:@9701.4]
  assign _T_9075 = offsetQ_5 < 4'he; // @[AxiLoadQueue.scala 131:33:@9702.4]
  assign _T_9078 = _T_9075 & _T_6368; // @[AxiLoadQueue.scala 131:41:@9704.4]
  assign _T_9080 = _T_9078 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9705.4]
  assign storesToCheck_5_14 = _T_2384 ? _T_9073 : _T_9080; // @[AxiLoadQueue.scala 130:10:@9706.4]
  assign _T_9086 = 4'hf <= offsetQ_5; // @[AxiLoadQueue.scala 130:81:@9709.4]
  assign storesToCheck_5_15 = _T_2384 ? _T_9086 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9715.4]
  assign storesToCheck_6_0 = _T_2414 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9757.4]
  assign _T_9136 = 4'h1 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9760.4]
  assign _T_9137 = _T_6138 & _T_9136; // @[AxiLoadQueue.scala 130:72:@9761.4]
  assign _T_9139 = offsetQ_6 < 4'h1; // @[AxiLoadQueue.scala 131:33:@9762.4]
  assign _T_9142 = _T_9139 & _T_6147; // @[AxiLoadQueue.scala 131:41:@9764.4]
  assign _T_9144 = _T_9142 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9765.4]
  assign storesToCheck_6_1 = _T_2414 ? _T_9137 : _T_9144; // @[AxiLoadQueue.scala 130:10:@9766.4]
  assign _T_9150 = 4'h2 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9769.4]
  assign _T_9151 = _T_6155 & _T_9150; // @[AxiLoadQueue.scala 130:72:@9770.4]
  assign _T_9153 = offsetQ_6 < 4'h2; // @[AxiLoadQueue.scala 131:33:@9771.4]
  assign _T_9156 = _T_9153 & _T_6164; // @[AxiLoadQueue.scala 131:41:@9773.4]
  assign _T_9158 = _T_9156 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9774.4]
  assign storesToCheck_6_2 = _T_2414 ? _T_9151 : _T_9158; // @[AxiLoadQueue.scala 130:10:@9775.4]
  assign _T_9164 = 4'h3 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9778.4]
  assign _T_9165 = _T_6172 & _T_9164; // @[AxiLoadQueue.scala 130:72:@9779.4]
  assign _T_9167 = offsetQ_6 < 4'h3; // @[AxiLoadQueue.scala 131:33:@9780.4]
  assign _T_9170 = _T_9167 & _T_6181; // @[AxiLoadQueue.scala 131:41:@9782.4]
  assign _T_9172 = _T_9170 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9783.4]
  assign storesToCheck_6_3 = _T_2414 ? _T_9165 : _T_9172; // @[AxiLoadQueue.scala 130:10:@9784.4]
  assign _T_9178 = 4'h4 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9787.4]
  assign _T_9179 = _T_6189 & _T_9178; // @[AxiLoadQueue.scala 130:72:@9788.4]
  assign _T_9181 = offsetQ_6 < 4'h4; // @[AxiLoadQueue.scala 131:33:@9789.4]
  assign _T_9184 = _T_9181 & _T_6198; // @[AxiLoadQueue.scala 131:41:@9791.4]
  assign _T_9186 = _T_9184 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9792.4]
  assign storesToCheck_6_4 = _T_2414 ? _T_9179 : _T_9186; // @[AxiLoadQueue.scala 130:10:@9793.4]
  assign _T_9192 = 4'h5 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9796.4]
  assign _T_9193 = _T_6206 & _T_9192; // @[AxiLoadQueue.scala 130:72:@9797.4]
  assign _T_9195 = offsetQ_6 < 4'h5; // @[AxiLoadQueue.scala 131:33:@9798.4]
  assign _T_9198 = _T_9195 & _T_6215; // @[AxiLoadQueue.scala 131:41:@9800.4]
  assign _T_9200 = _T_9198 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9801.4]
  assign storesToCheck_6_5 = _T_2414 ? _T_9193 : _T_9200; // @[AxiLoadQueue.scala 130:10:@9802.4]
  assign _T_9206 = 4'h6 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9805.4]
  assign _T_9207 = _T_6223 & _T_9206; // @[AxiLoadQueue.scala 130:72:@9806.4]
  assign _T_9209 = offsetQ_6 < 4'h6; // @[AxiLoadQueue.scala 131:33:@9807.4]
  assign _T_9212 = _T_9209 & _T_6232; // @[AxiLoadQueue.scala 131:41:@9809.4]
  assign _T_9214 = _T_9212 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9810.4]
  assign storesToCheck_6_6 = _T_2414 ? _T_9207 : _T_9214; // @[AxiLoadQueue.scala 130:10:@9811.4]
  assign _T_9220 = 4'h7 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9814.4]
  assign _T_9221 = _T_6240 & _T_9220; // @[AxiLoadQueue.scala 130:72:@9815.4]
  assign _T_9223 = offsetQ_6 < 4'h7; // @[AxiLoadQueue.scala 131:33:@9816.4]
  assign _T_9226 = _T_9223 & _T_6249; // @[AxiLoadQueue.scala 131:41:@9818.4]
  assign _T_9228 = _T_9226 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9819.4]
  assign storesToCheck_6_7 = _T_2414 ? _T_9221 : _T_9228; // @[AxiLoadQueue.scala 130:10:@9820.4]
  assign _T_9234 = 4'h8 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9823.4]
  assign _T_9235 = _T_6257 & _T_9234; // @[AxiLoadQueue.scala 130:72:@9824.4]
  assign _T_9237 = offsetQ_6 < 4'h8; // @[AxiLoadQueue.scala 131:33:@9825.4]
  assign _T_9240 = _T_9237 & _T_6266; // @[AxiLoadQueue.scala 131:41:@9827.4]
  assign _T_9242 = _T_9240 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9828.4]
  assign storesToCheck_6_8 = _T_2414 ? _T_9235 : _T_9242; // @[AxiLoadQueue.scala 130:10:@9829.4]
  assign _T_9248 = 4'h9 <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9832.4]
  assign _T_9249 = _T_6274 & _T_9248; // @[AxiLoadQueue.scala 130:72:@9833.4]
  assign _T_9251 = offsetQ_6 < 4'h9; // @[AxiLoadQueue.scala 131:33:@9834.4]
  assign _T_9254 = _T_9251 & _T_6283; // @[AxiLoadQueue.scala 131:41:@9836.4]
  assign _T_9256 = _T_9254 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9837.4]
  assign storesToCheck_6_9 = _T_2414 ? _T_9249 : _T_9256; // @[AxiLoadQueue.scala 130:10:@9838.4]
  assign _T_9262 = 4'ha <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9841.4]
  assign _T_9263 = _T_6291 & _T_9262; // @[AxiLoadQueue.scala 130:72:@9842.4]
  assign _T_9265 = offsetQ_6 < 4'ha; // @[AxiLoadQueue.scala 131:33:@9843.4]
  assign _T_9268 = _T_9265 & _T_6300; // @[AxiLoadQueue.scala 131:41:@9845.4]
  assign _T_9270 = _T_9268 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9846.4]
  assign storesToCheck_6_10 = _T_2414 ? _T_9263 : _T_9270; // @[AxiLoadQueue.scala 130:10:@9847.4]
  assign _T_9276 = 4'hb <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9850.4]
  assign _T_9277 = _T_6308 & _T_9276; // @[AxiLoadQueue.scala 130:72:@9851.4]
  assign _T_9279 = offsetQ_6 < 4'hb; // @[AxiLoadQueue.scala 131:33:@9852.4]
  assign _T_9282 = _T_9279 & _T_6317; // @[AxiLoadQueue.scala 131:41:@9854.4]
  assign _T_9284 = _T_9282 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9855.4]
  assign storesToCheck_6_11 = _T_2414 ? _T_9277 : _T_9284; // @[AxiLoadQueue.scala 130:10:@9856.4]
  assign _T_9290 = 4'hc <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9859.4]
  assign _T_9291 = _T_6325 & _T_9290; // @[AxiLoadQueue.scala 130:72:@9860.4]
  assign _T_9293 = offsetQ_6 < 4'hc; // @[AxiLoadQueue.scala 131:33:@9861.4]
  assign _T_9296 = _T_9293 & _T_6334; // @[AxiLoadQueue.scala 131:41:@9863.4]
  assign _T_9298 = _T_9296 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9864.4]
  assign storesToCheck_6_12 = _T_2414 ? _T_9291 : _T_9298; // @[AxiLoadQueue.scala 130:10:@9865.4]
  assign _T_9304 = 4'hd <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9868.4]
  assign _T_9305 = _T_6342 & _T_9304; // @[AxiLoadQueue.scala 130:72:@9869.4]
  assign _T_9307 = offsetQ_6 < 4'hd; // @[AxiLoadQueue.scala 131:33:@9870.4]
  assign _T_9310 = _T_9307 & _T_6351; // @[AxiLoadQueue.scala 131:41:@9872.4]
  assign _T_9312 = _T_9310 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9873.4]
  assign storesToCheck_6_13 = _T_2414 ? _T_9305 : _T_9312; // @[AxiLoadQueue.scala 130:10:@9874.4]
  assign _T_9318 = 4'he <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9877.4]
  assign _T_9319 = _T_6359 & _T_9318; // @[AxiLoadQueue.scala 130:72:@9878.4]
  assign _T_9321 = offsetQ_6 < 4'he; // @[AxiLoadQueue.scala 131:33:@9879.4]
  assign _T_9324 = _T_9321 & _T_6368; // @[AxiLoadQueue.scala 131:41:@9881.4]
  assign _T_9326 = _T_9324 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9882.4]
  assign storesToCheck_6_14 = _T_2414 ? _T_9319 : _T_9326; // @[AxiLoadQueue.scala 130:10:@9883.4]
  assign _T_9332 = 4'hf <= offsetQ_6; // @[AxiLoadQueue.scala 130:81:@9886.4]
  assign storesToCheck_6_15 = _T_2414 ? _T_9332 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9892.4]
  assign storesToCheck_7_0 = _T_2444 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@9934.4]
  assign _T_9382 = 4'h1 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@9937.4]
  assign _T_9383 = _T_6138 & _T_9382; // @[AxiLoadQueue.scala 130:72:@9938.4]
  assign _T_9385 = offsetQ_7 < 4'h1; // @[AxiLoadQueue.scala 131:33:@9939.4]
  assign _T_9388 = _T_9385 & _T_6147; // @[AxiLoadQueue.scala 131:41:@9941.4]
  assign _T_9390 = _T_9388 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9942.4]
  assign storesToCheck_7_1 = _T_2444 ? _T_9383 : _T_9390; // @[AxiLoadQueue.scala 130:10:@9943.4]
  assign _T_9396 = 4'h2 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@9946.4]
  assign _T_9397 = _T_6155 & _T_9396; // @[AxiLoadQueue.scala 130:72:@9947.4]
  assign _T_9399 = offsetQ_7 < 4'h2; // @[AxiLoadQueue.scala 131:33:@9948.4]
  assign _T_9402 = _T_9399 & _T_6164; // @[AxiLoadQueue.scala 131:41:@9950.4]
  assign _T_9404 = _T_9402 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9951.4]
  assign storesToCheck_7_2 = _T_2444 ? _T_9397 : _T_9404; // @[AxiLoadQueue.scala 130:10:@9952.4]
  assign _T_9410 = 4'h3 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@9955.4]
  assign _T_9411 = _T_6172 & _T_9410; // @[AxiLoadQueue.scala 130:72:@9956.4]
  assign _T_9413 = offsetQ_7 < 4'h3; // @[AxiLoadQueue.scala 131:33:@9957.4]
  assign _T_9416 = _T_9413 & _T_6181; // @[AxiLoadQueue.scala 131:41:@9959.4]
  assign _T_9418 = _T_9416 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9960.4]
  assign storesToCheck_7_3 = _T_2444 ? _T_9411 : _T_9418; // @[AxiLoadQueue.scala 130:10:@9961.4]
  assign _T_9424 = 4'h4 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@9964.4]
  assign _T_9425 = _T_6189 & _T_9424; // @[AxiLoadQueue.scala 130:72:@9965.4]
  assign _T_9427 = offsetQ_7 < 4'h4; // @[AxiLoadQueue.scala 131:33:@9966.4]
  assign _T_9430 = _T_9427 & _T_6198; // @[AxiLoadQueue.scala 131:41:@9968.4]
  assign _T_9432 = _T_9430 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9969.4]
  assign storesToCheck_7_4 = _T_2444 ? _T_9425 : _T_9432; // @[AxiLoadQueue.scala 130:10:@9970.4]
  assign _T_9438 = 4'h5 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@9973.4]
  assign _T_9439 = _T_6206 & _T_9438; // @[AxiLoadQueue.scala 130:72:@9974.4]
  assign _T_9441 = offsetQ_7 < 4'h5; // @[AxiLoadQueue.scala 131:33:@9975.4]
  assign _T_9444 = _T_9441 & _T_6215; // @[AxiLoadQueue.scala 131:41:@9977.4]
  assign _T_9446 = _T_9444 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9978.4]
  assign storesToCheck_7_5 = _T_2444 ? _T_9439 : _T_9446; // @[AxiLoadQueue.scala 130:10:@9979.4]
  assign _T_9452 = 4'h6 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@9982.4]
  assign _T_9453 = _T_6223 & _T_9452; // @[AxiLoadQueue.scala 130:72:@9983.4]
  assign _T_9455 = offsetQ_7 < 4'h6; // @[AxiLoadQueue.scala 131:33:@9984.4]
  assign _T_9458 = _T_9455 & _T_6232; // @[AxiLoadQueue.scala 131:41:@9986.4]
  assign _T_9460 = _T_9458 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9987.4]
  assign storesToCheck_7_6 = _T_2444 ? _T_9453 : _T_9460; // @[AxiLoadQueue.scala 130:10:@9988.4]
  assign _T_9466 = 4'h7 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@9991.4]
  assign _T_9467 = _T_6240 & _T_9466; // @[AxiLoadQueue.scala 130:72:@9992.4]
  assign _T_9469 = offsetQ_7 < 4'h7; // @[AxiLoadQueue.scala 131:33:@9993.4]
  assign _T_9472 = _T_9469 & _T_6249; // @[AxiLoadQueue.scala 131:41:@9995.4]
  assign _T_9474 = _T_9472 == 1'h0; // @[AxiLoadQueue.scala 131:9:@9996.4]
  assign storesToCheck_7_7 = _T_2444 ? _T_9467 : _T_9474; // @[AxiLoadQueue.scala 130:10:@9997.4]
  assign _T_9480 = 4'h8 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10000.4]
  assign _T_9481 = _T_6257 & _T_9480; // @[AxiLoadQueue.scala 130:72:@10001.4]
  assign _T_9483 = offsetQ_7 < 4'h8; // @[AxiLoadQueue.scala 131:33:@10002.4]
  assign _T_9486 = _T_9483 & _T_6266; // @[AxiLoadQueue.scala 131:41:@10004.4]
  assign _T_9488 = _T_9486 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10005.4]
  assign storesToCheck_7_8 = _T_2444 ? _T_9481 : _T_9488; // @[AxiLoadQueue.scala 130:10:@10006.4]
  assign _T_9494 = 4'h9 <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10009.4]
  assign _T_9495 = _T_6274 & _T_9494; // @[AxiLoadQueue.scala 130:72:@10010.4]
  assign _T_9497 = offsetQ_7 < 4'h9; // @[AxiLoadQueue.scala 131:33:@10011.4]
  assign _T_9500 = _T_9497 & _T_6283; // @[AxiLoadQueue.scala 131:41:@10013.4]
  assign _T_9502 = _T_9500 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10014.4]
  assign storesToCheck_7_9 = _T_2444 ? _T_9495 : _T_9502; // @[AxiLoadQueue.scala 130:10:@10015.4]
  assign _T_9508 = 4'ha <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10018.4]
  assign _T_9509 = _T_6291 & _T_9508; // @[AxiLoadQueue.scala 130:72:@10019.4]
  assign _T_9511 = offsetQ_7 < 4'ha; // @[AxiLoadQueue.scala 131:33:@10020.4]
  assign _T_9514 = _T_9511 & _T_6300; // @[AxiLoadQueue.scala 131:41:@10022.4]
  assign _T_9516 = _T_9514 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10023.4]
  assign storesToCheck_7_10 = _T_2444 ? _T_9509 : _T_9516; // @[AxiLoadQueue.scala 130:10:@10024.4]
  assign _T_9522 = 4'hb <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10027.4]
  assign _T_9523 = _T_6308 & _T_9522; // @[AxiLoadQueue.scala 130:72:@10028.4]
  assign _T_9525 = offsetQ_7 < 4'hb; // @[AxiLoadQueue.scala 131:33:@10029.4]
  assign _T_9528 = _T_9525 & _T_6317; // @[AxiLoadQueue.scala 131:41:@10031.4]
  assign _T_9530 = _T_9528 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10032.4]
  assign storesToCheck_7_11 = _T_2444 ? _T_9523 : _T_9530; // @[AxiLoadQueue.scala 130:10:@10033.4]
  assign _T_9536 = 4'hc <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10036.4]
  assign _T_9537 = _T_6325 & _T_9536; // @[AxiLoadQueue.scala 130:72:@10037.4]
  assign _T_9539 = offsetQ_7 < 4'hc; // @[AxiLoadQueue.scala 131:33:@10038.4]
  assign _T_9542 = _T_9539 & _T_6334; // @[AxiLoadQueue.scala 131:41:@10040.4]
  assign _T_9544 = _T_9542 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10041.4]
  assign storesToCheck_7_12 = _T_2444 ? _T_9537 : _T_9544; // @[AxiLoadQueue.scala 130:10:@10042.4]
  assign _T_9550 = 4'hd <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10045.4]
  assign _T_9551 = _T_6342 & _T_9550; // @[AxiLoadQueue.scala 130:72:@10046.4]
  assign _T_9553 = offsetQ_7 < 4'hd; // @[AxiLoadQueue.scala 131:33:@10047.4]
  assign _T_9556 = _T_9553 & _T_6351; // @[AxiLoadQueue.scala 131:41:@10049.4]
  assign _T_9558 = _T_9556 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10050.4]
  assign storesToCheck_7_13 = _T_2444 ? _T_9551 : _T_9558; // @[AxiLoadQueue.scala 130:10:@10051.4]
  assign _T_9564 = 4'he <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10054.4]
  assign _T_9565 = _T_6359 & _T_9564; // @[AxiLoadQueue.scala 130:72:@10055.4]
  assign _T_9567 = offsetQ_7 < 4'he; // @[AxiLoadQueue.scala 131:33:@10056.4]
  assign _T_9570 = _T_9567 & _T_6368; // @[AxiLoadQueue.scala 131:41:@10058.4]
  assign _T_9572 = _T_9570 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10059.4]
  assign storesToCheck_7_14 = _T_2444 ? _T_9565 : _T_9572; // @[AxiLoadQueue.scala 130:10:@10060.4]
  assign _T_9578 = 4'hf <= offsetQ_7; // @[AxiLoadQueue.scala 130:81:@10063.4]
  assign storesToCheck_7_15 = _T_2444 ? _T_9578 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10069.4]
  assign storesToCheck_8_0 = _T_2474 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10111.4]
  assign _T_9628 = 4'h1 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10114.4]
  assign _T_9629 = _T_6138 & _T_9628; // @[AxiLoadQueue.scala 130:72:@10115.4]
  assign _T_9631 = offsetQ_8 < 4'h1; // @[AxiLoadQueue.scala 131:33:@10116.4]
  assign _T_9634 = _T_9631 & _T_6147; // @[AxiLoadQueue.scala 131:41:@10118.4]
  assign _T_9636 = _T_9634 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10119.4]
  assign storesToCheck_8_1 = _T_2474 ? _T_9629 : _T_9636; // @[AxiLoadQueue.scala 130:10:@10120.4]
  assign _T_9642 = 4'h2 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10123.4]
  assign _T_9643 = _T_6155 & _T_9642; // @[AxiLoadQueue.scala 130:72:@10124.4]
  assign _T_9645 = offsetQ_8 < 4'h2; // @[AxiLoadQueue.scala 131:33:@10125.4]
  assign _T_9648 = _T_9645 & _T_6164; // @[AxiLoadQueue.scala 131:41:@10127.4]
  assign _T_9650 = _T_9648 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10128.4]
  assign storesToCheck_8_2 = _T_2474 ? _T_9643 : _T_9650; // @[AxiLoadQueue.scala 130:10:@10129.4]
  assign _T_9656 = 4'h3 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10132.4]
  assign _T_9657 = _T_6172 & _T_9656; // @[AxiLoadQueue.scala 130:72:@10133.4]
  assign _T_9659 = offsetQ_8 < 4'h3; // @[AxiLoadQueue.scala 131:33:@10134.4]
  assign _T_9662 = _T_9659 & _T_6181; // @[AxiLoadQueue.scala 131:41:@10136.4]
  assign _T_9664 = _T_9662 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10137.4]
  assign storesToCheck_8_3 = _T_2474 ? _T_9657 : _T_9664; // @[AxiLoadQueue.scala 130:10:@10138.4]
  assign _T_9670 = 4'h4 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10141.4]
  assign _T_9671 = _T_6189 & _T_9670; // @[AxiLoadQueue.scala 130:72:@10142.4]
  assign _T_9673 = offsetQ_8 < 4'h4; // @[AxiLoadQueue.scala 131:33:@10143.4]
  assign _T_9676 = _T_9673 & _T_6198; // @[AxiLoadQueue.scala 131:41:@10145.4]
  assign _T_9678 = _T_9676 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10146.4]
  assign storesToCheck_8_4 = _T_2474 ? _T_9671 : _T_9678; // @[AxiLoadQueue.scala 130:10:@10147.4]
  assign _T_9684 = 4'h5 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10150.4]
  assign _T_9685 = _T_6206 & _T_9684; // @[AxiLoadQueue.scala 130:72:@10151.4]
  assign _T_9687 = offsetQ_8 < 4'h5; // @[AxiLoadQueue.scala 131:33:@10152.4]
  assign _T_9690 = _T_9687 & _T_6215; // @[AxiLoadQueue.scala 131:41:@10154.4]
  assign _T_9692 = _T_9690 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10155.4]
  assign storesToCheck_8_5 = _T_2474 ? _T_9685 : _T_9692; // @[AxiLoadQueue.scala 130:10:@10156.4]
  assign _T_9698 = 4'h6 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10159.4]
  assign _T_9699 = _T_6223 & _T_9698; // @[AxiLoadQueue.scala 130:72:@10160.4]
  assign _T_9701 = offsetQ_8 < 4'h6; // @[AxiLoadQueue.scala 131:33:@10161.4]
  assign _T_9704 = _T_9701 & _T_6232; // @[AxiLoadQueue.scala 131:41:@10163.4]
  assign _T_9706 = _T_9704 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10164.4]
  assign storesToCheck_8_6 = _T_2474 ? _T_9699 : _T_9706; // @[AxiLoadQueue.scala 130:10:@10165.4]
  assign _T_9712 = 4'h7 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10168.4]
  assign _T_9713 = _T_6240 & _T_9712; // @[AxiLoadQueue.scala 130:72:@10169.4]
  assign _T_9715 = offsetQ_8 < 4'h7; // @[AxiLoadQueue.scala 131:33:@10170.4]
  assign _T_9718 = _T_9715 & _T_6249; // @[AxiLoadQueue.scala 131:41:@10172.4]
  assign _T_9720 = _T_9718 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10173.4]
  assign storesToCheck_8_7 = _T_2474 ? _T_9713 : _T_9720; // @[AxiLoadQueue.scala 130:10:@10174.4]
  assign _T_9726 = 4'h8 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10177.4]
  assign _T_9727 = _T_6257 & _T_9726; // @[AxiLoadQueue.scala 130:72:@10178.4]
  assign _T_9729 = offsetQ_8 < 4'h8; // @[AxiLoadQueue.scala 131:33:@10179.4]
  assign _T_9732 = _T_9729 & _T_6266; // @[AxiLoadQueue.scala 131:41:@10181.4]
  assign _T_9734 = _T_9732 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10182.4]
  assign storesToCheck_8_8 = _T_2474 ? _T_9727 : _T_9734; // @[AxiLoadQueue.scala 130:10:@10183.4]
  assign _T_9740 = 4'h9 <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10186.4]
  assign _T_9741 = _T_6274 & _T_9740; // @[AxiLoadQueue.scala 130:72:@10187.4]
  assign _T_9743 = offsetQ_8 < 4'h9; // @[AxiLoadQueue.scala 131:33:@10188.4]
  assign _T_9746 = _T_9743 & _T_6283; // @[AxiLoadQueue.scala 131:41:@10190.4]
  assign _T_9748 = _T_9746 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10191.4]
  assign storesToCheck_8_9 = _T_2474 ? _T_9741 : _T_9748; // @[AxiLoadQueue.scala 130:10:@10192.4]
  assign _T_9754 = 4'ha <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10195.4]
  assign _T_9755 = _T_6291 & _T_9754; // @[AxiLoadQueue.scala 130:72:@10196.4]
  assign _T_9757 = offsetQ_8 < 4'ha; // @[AxiLoadQueue.scala 131:33:@10197.4]
  assign _T_9760 = _T_9757 & _T_6300; // @[AxiLoadQueue.scala 131:41:@10199.4]
  assign _T_9762 = _T_9760 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10200.4]
  assign storesToCheck_8_10 = _T_2474 ? _T_9755 : _T_9762; // @[AxiLoadQueue.scala 130:10:@10201.4]
  assign _T_9768 = 4'hb <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10204.4]
  assign _T_9769 = _T_6308 & _T_9768; // @[AxiLoadQueue.scala 130:72:@10205.4]
  assign _T_9771 = offsetQ_8 < 4'hb; // @[AxiLoadQueue.scala 131:33:@10206.4]
  assign _T_9774 = _T_9771 & _T_6317; // @[AxiLoadQueue.scala 131:41:@10208.4]
  assign _T_9776 = _T_9774 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10209.4]
  assign storesToCheck_8_11 = _T_2474 ? _T_9769 : _T_9776; // @[AxiLoadQueue.scala 130:10:@10210.4]
  assign _T_9782 = 4'hc <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10213.4]
  assign _T_9783 = _T_6325 & _T_9782; // @[AxiLoadQueue.scala 130:72:@10214.4]
  assign _T_9785 = offsetQ_8 < 4'hc; // @[AxiLoadQueue.scala 131:33:@10215.4]
  assign _T_9788 = _T_9785 & _T_6334; // @[AxiLoadQueue.scala 131:41:@10217.4]
  assign _T_9790 = _T_9788 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10218.4]
  assign storesToCheck_8_12 = _T_2474 ? _T_9783 : _T_9790; // @[AxiLoadQueue.scala 130:10:@10219.4]
  assign _T_9796 = 4'hd <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10222.4]
  assign _T_9797 = _T_6342 & _T_9796; // @[AxiLoadQueue.scala 130:72:@10223.4]
  assign _T_9799 = offsetQ_8 < 4'hd; // @[AxiLoadQueue.scala 131:33:@10224.4]
  assign _T_9802 = _T_9799 & _T_6351; // @[AxiLoadQueue.scala 131:41:@10226.4]
  assign _T_9804 = _T_9802 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10227.4]
  assign storesToCheck_8_13 = _T_2474 ? _T_9797 : _T_9804; // @[AxiLoadQueue.scala 130:10:@10228.4]
  assign _T_9810 = 4'he <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10231.4]
  assign _T_9811 = _T_6359 & _T_9810; // @[AxiLoadQueue.scala 130:72:@10232.4]
  assign _T_9813 = offsetQ_8 < 4'he; // @[AxiLoadQueue.scala 131:33:@10233.4]
  assign _T_9816 = _T_9813 & _T_6368; // @[AxiLoadQueue.scala 131:41:@10235.4]
  assign _T_9818 = _T_9816 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10236.4]
  assign storesToCheck_8_14 = _T_2474 ? _T_9811 : _T_9818; // @[AxiLoadQueue.scala 130:10:@10237.4]
  assign _T_9824 = 4'hf <= offsetQ_8; // @[AxiLoadQueue.scala 130:81:@10240.4]
  assign storesToCheck_8_15 = _T_2474 ? _T_9824 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10246.4]
  assign storesToCheck_9_0 = _T_2504 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10288.4]
  assign _T_9874 = 4'h1 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10291.4]
  assign _T_9875 = _T_6138 & _T_9874; // @[AxiLoadQueue.scala 130:72:@10292.4]
  assign _T_9877 = offsetQ_9 < 4'h1; // @[AxiLoadQueue.scala 131:33:@10293.4]
  assign _T_9880 = _T_9877 & _T_6147; // @[AxiLoadQueue.scala 131:41:@10295.4]
  assign _T_9882 = _T_9880 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10296.4]
  assign storesToCheck_9_1 = _T_2504 ? _T_9875 : _T_9882; // @[AxiLoadQueue.scala 130:10:@10297.4]
  assign _T_9888 = 4'h2 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10300.4]
  assign _T_9889 = _T_6155 & _T_9888; // @[AxiLoadQueue.scala 130:72:@10301.4]
  assign _T_9891 = offsetQ_9 < 4'h2; // @[AxiLoadQueue.scala 131:33:@10302.4]
  assign _T_9894 = _T_9891 & _T_6164; // @[AxiLoadQueue.scala 131:41:@10304.4]
  assign _T_9896 = _T_9894 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10305.4]
  assign storesToCheck_9_2 = _T_2504 ? _T_9889 : _T_9896; // @[AxiLoadQueue.scala 130:10:@10306.4]
  assign _T_9902 = 4'h3 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10309.4]
  assign _T_9903 = _T_6172 & _T_9902; // @[AxiLoadQueue.scala 130:72:@10310.4]
  assign _T_9905 = offsetQ_9 < 4'h3; // @[AxiLoadQueue.scala 131:33:@10311.4]
  assign _T_9908 = _T_9905 & _T_6181; // @[AxiLoadQueue.scala 131:41:@10313.4]
  assign _T_9910 = _T_9908 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10314.4]
  assign storesToCheck_9_3 = _T_2504 ? _T_9903 : _T_9910; // @[AxiLoadQueue.scala 130:10:@10315.4]
  assign _T_9916 = 4'h4 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10318.4]
  assign _T_9917 = _T_6189 & _T_9916; // @[AxiLoadQueue.scala 130:72:@10319.4]
  assign _T_9919 = offsetQ_9 < 4'h4; // @[AxiLoadQueue.scala 131:33:@10320.4]
  assign _T_9922 = _T_9919 & _T_6198; // @[AxiLoadQueue.scala 131:41:@10322.4]
  assign _T_9924 = _T_9922 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10323.4]
  assign storesToCheck_9_4 = _T_2504 ? _T_9917 : _T_9924; // @[AxiLoadQueue.scala 130:10:@10324.4]
  assign _T_9930 = 4'h5 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10327.4]
  assign _T_9931 = _T_6206 & _T_9930; // @[AxiLoadQueue.scala 130:72:@10328.4]
  assign _T_9933 = offsetQ_9 < 4'h5; // @[AxiLoadQueue.scala 131:33:@10329.4]
  assign _T_9936 = _T_9933 & _T_6215; // @[AxiLoadQueue.scala 131:41:@10331.4]
  assign _T_9938 = _T_9936 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10332.4]
  assign storesToCheck_9_5 = _T_2504 ? _T_9931 : _T_9938; // @[AxiLoadQueue.scala 130:10:@10333.4]
  assign _T_9944 = 4'h6 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10336.4]
  assign _T_9945 = _T_6223 & _T_9944; // @[AxiLoadQueue.scala 130:72:@10337.4]
  assign _T_9947 = offsetQ_9 < 4'h6; // @[AxiLoadQueue.scala 131:33:@10338.4]
  assign _T_9950 = _T_9947 & _T_6232; // @[AxiLoadQueue.scala 131:41:@10340.4]
  assign _T_9952 = _T_9950 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10341.4]
  assign storesToCheck_9_6 = _T_2504 ? _T_9945 : _T_9952; // @[AxiLoadQueue.scala 130:10:@10342.4]
  assign _T_9958 = 4'h7 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10345.4]
  assign _T_9959 = _T_6240 & _T_9958; // @[AxiLoadQueue.scala 130:72:@10346.4]
  assign _T_9961 = offsetQ_9 < 4'h7; // @[AxiLoadQueue.scala 131:33:@10347.4]
  assign _T_9964 = _T_9961 & _T_6249; // @[AxiLoadQueue.scala 131:41:@10349.4]
  assign _T_9966 = _T_9964 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10350.4]
  assign storesToCheck_9_7 = _T_2504 ? _T_9959 : _T_9966; // @[AxiLoadQueue.scala 130:10:@10351.4]
  assign _T_9972 = 4'h8 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10354.4]
  assign _T_9973 = _T_6257 & _T_9972; // @[AxiLoadQueue.scala 130:72:@10355.4]
  assign _T_9975 = offsetQ_9 < 4'h8; // @[AxiLoadQueue.scala 131:33:@10356.4]
  assign _T_9978 = _T_9975 & _T_6266; // @[AxiLoadQueue.scala 131:41:@10358.4]
  assign _T_9980 = _T_9978 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10359.4]
  assign storesToCheck_9_8 = _T_2504 ? _T_9973 : _T_9980; // @[AxiLoadQueue.scala 130:10:@10360.4]
  assign _T_9986 = 4'h9 <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10363.4]
  assign _T_9987 = _T_6274 & _T_9986; // @[AxiLoadQueue.scala 130:72:@10364.4]
  assign _T_9989 = offsetQ_9 < 4'h9; // @[AxiLoadQueue.scala 131:33:@10365.4]
  assign _T_9992 = _T_9989 & _T_6283; // @[AxiLoadQueue.scala 131:41:@10367.4]
  assign _T_9994 = _T_9992 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10368.4]
  assign storesToCheck_9_9 = _T_2504 ? _T_9987 : _T_9994; // @[AxiLoadQueue.scala 130:10:@10369.4]
  assign _T_10000 = 4'ha <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10372.4]
  assign _T_10001 = _T_6291 & _T_10000; // @[AxiLoadQueue.scala 130:72:@10373.4]
  assign _T_10003 = offsetQ_9 < 4'ha; // @[AxiLoadQueue.scala 131:33:@10374.4]
  assign _T_10006 = _T_10003 & _T_6300; // @[AxiLoadQueue.scala 131:41:@10376.4]
  assign _T_10008 = _T_10006 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10377.4]
  assign storesToCheck_9_10 = _T_2504 ? _T_10001 : _T_10008; // @[AxiLoadQueue.scala 130:10:@10378.4]
  assign _T_10014 = 4'hb <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10381.4]
  assign _T_10015 = _T_6308 & _T_10014; // @[AxiLoadQueue.scala 130:72:@10382.4]
  assign _T_10017 = offsetQ_9 < 4'hb; // @[AxiLoadQueue.scala 131:33:@10383.4]
  assign _T_10020 = _T_10017 & _T_6317; // @[AxiLoadQueue.scala 131:41:@10385.4]
  assign _T_10022 = _T_10020 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10386.4]
  assign storesToCheck_9_11 = _T_2504 ? _T_10015 : _T_10022; // @[AxiLoadQueue.scala 130:10:@10387.4]
  assign _T_10028 = 4'hc <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10390.4]
  assign _T_10029 = _T_6325 & _T_10028; // @[AxiLoadQueue.scala 130:72:@10391.4]
  assign _T_10031 = offsetQ_9 < 4'hc; // @[AxiLoadQueue.scala 131:33:@10392.4]
  assign _T_10034 = _T_10031 & _T_6334; // @[AxiLoadQueue.scala 131:41:@10394.4]
  assign _T_10036 = _T_10034 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10395.4]
  assign storesToCheck_9_12 = _T_2504 ? _T_10029 : _T_10036; // @[AxiLoadQueue.scala 130:10:@10396.4]
  assign _T_10042 = 4'hd <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10399.4]
  assign _T_10043 = _T_6342 & _T_10042; // @[AxiLoadQueue.scala 130:72:@10400.4]
  assign _T_10045 = offsetQ_9 < 4'hd; // @[AxiLoadQueue.scala 131:33:@10401.4]
  assign _T_10048 = _T_10045 & _T_6351; // @[AxiLoadQueue.scala 131:41:@10403.4]
  assign _T_10050 = _T_10048 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10404.4]
  assign storesToCheck_9_13 = _T_2504 ? _T_10043 : _T_10050; // @[AxiLoadQueue.scala 130:10:@10405.4]
  assign _T_10056 = 4'he <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10408.4]
  assign _T_10057 = _T_6359 & _T_10056; // @[AxiLoadQueue.scala 130:72:@10409.4]
  assign _T_10059 = offsetQ_9 < 4'he; // @[AxiLoadQueue.scala 131:33:@10410.4]
  assign _T_10062 = _T_10059 & _T_6368; // @[AxiLoadQueue.scala 131:41:@10412.4]
  assign _T_10064 = _T_10062 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10413.4]
  assign storesToCheck_9_14 = _T_2504 ? _T_10057 : _T_10064; // @[AxiLoadQueue.scala 130:10:@10414.4]
  assign _T_10070 = 4'hf <= offsetQ_9; // @[AxiLoadQueue.scala 130:81:@10417.4]
  assign storesToCheck_9_15 = _T_2504 ? _T_10070 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10423.4]
  assign storesToCheck_10_0 = _T_2534 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10465.4]
  assign _T_10120 = 4'h1 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10468.4]
  assign _T_10121 = _T_6138 & _T_10120; // @[AxiLoadQueue.scala 130:72:@10469.4]
  assign _T_10123 = offsetQ_10 < 4'h1; // @[AxiLoadQueue.scala 131:33:@10470.4]
  assign _T_10126 = _T_10123 & _T_6147; // @[AxiLoadQueue.scala 131:41:@10472.4]
  assign _T_10128 = _T_10126 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10473.4]
  assign storesToCheck_10_1 = _T_2534 ? _T_10121 : _T_10128; // @[AxiLoadQueue.scala 130:10:@10474.4]
  assign _T_10134 = 4'h2 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10477.4]
  assign _T_10135 = _T_6155 & _T_10134; // @[AxiLoadQueue.scala 130:72:@10478.4]
  assign _T_10137 = offsetQ_10 < 4'h2; // @[AxiLoadQueue.scala 131:33:@10479.4]
  assign _T_10140 = _T_10137 & _T_6164; // @[AxiLoadQueue.scala 131:41:@10481.4]
  assign _T_10142 = _T_10140 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10482.4]
  assign storesToCheck_10_2 = _T_2534 ? _T_10135 : _T_10142; // @[AxiLoadQueue.scala 130:10:@10483.4]
  assign _T_10148 = 4'h3 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10486.4]
  assign _T_10149 = _T_6172 & _T_10148; // @[AxiLoadQueue.scala 130:72:@10487.4]
  assign _T_10151 = offsetQ_10 < 4'h3; // @[AxiLoadQueue.scala 131:33:@10488.4]
  assign _T_10154 = _T_10151 & _T_6181; // @[AxiLoadQueue.scala 131:41:@10490.4]
  assign _T_10156 = _T_10154 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10491.4]
  assign storesToCheck_10_3 = _T_2534 ? _T_10149 : _T_10156; // @[AxiLoadQueue.scala 130:10:@10492.4]
  assign _T_10162 = 4'h4 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10495.4]
  assign _T_10163 = _T_6189 & _T_10162; // @[AxiLoadQueue.scala 130:72:@10496.4]
  assign _T_10165 = offsetQ_10 < 4'h4; // @[AxiLoadQueue.scala 131:33:@10497.4]
  assign _T_10168 = _T_10165 & _T_6198; // @[AxiLoadQueue.scala 131:41:@10499.4]
  assign _T_10170 = _T_10168 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10500.4]
  assign storesToCheck_10_4 = _T_2534 ? _T_10163 : _T_10170; // @[AxiLoadQueue.scala 130:10:@10501.4]
  assign _T_10176 = 4'h5 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10504.4]
  assign _T_10177 = _T_6206 & _T_10176; // @[AxiLoadQueue.scala 130:72:@10505.4]
  assign _T_10179 = offsetQ_10 < 4'h5; // @[AxiLoadQueue.scala 131:33:@10506.4]
  assign _T_10182 = _T_10179 & _T_6215; // @[AxiLoadQueue.scala 131:41:@10508.4]
  assign _T_10184 = _T_10182 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10509.4]
  assign storesToCheck_10_5 = _T_2534 ? _T_10177 : _T_10184; // @[AxiLoadQueue.scala 130:10:@10510.4]
  assign _T_10190 = 4'h6 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10513.4]
  assign _T_10191 = _T_6223 & _T_10190; // @[AxiLoadQueue.scala 130:72:@10514.4]
  assign _T_10193 = offsetQ_10 < 4'h6; // @[AxiLoadQueue.scala 131:33:@10515.4]
  assign _T_10196 = _T_10193 & _T_6232; // @[AxiLoadQueue.scala 131:41:@10517.4]
  assign _T_10198 = _T_10196 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10518.4]
  assign storesToCheck_10_6 = _T_2534 ? _T_10191 : _T_10198; // @[AxiLoadQueue.scala 130:10:@10519.4]
  assign _T_10204 = 4'h7 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10522.4]
  assign _T_10205 = _T_6240 & _T_10204; // @[AxiLoadQueue.scala 130:72:@10523.4]
  assign _T_10207 = offsetQ_10 < 4'h7; // @[AxiLoadQueue.scala 131:33:@10524.4]
  assign _T_10210 = _T_10207 & _T_6249; // @[AxiLoadQueue.scala 131:41:@10526.4]
  assign _T_10212 = _T_10210 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10527.4]
  assign storesToCheck_10_7 = _T_2534 ? _T_10205 : _T_10212; // @[AxiLoadQueue.scala 130:10:@10528.4]
  assign _T_10218 = 4'h8 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10531.4]
  assign _T_10219 = _T_6257 & _T_10218; // @[AxiLoadQueue.scala 130:72:@10532.4]
  assign _T_10221 = offsetQ_10 < 4'h8; // @[AxiLoadQueue.scala 131:33:@10533.4]
  assign _T_10224 = _T_10221 & _T_6266; // @[AxiLoadQueue.scala 131:41:@10535.4]
  assign _T_10226 = _T_10224 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10536.4]
  assign storesToCheck_10_8 = _T_2534 ? _T_10219 : _T_10226; // @[AxiLoadQueue.scala 130:10:@10537.4]
  assign _T_10232 = 4'h9 <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10540.4]
  assign _T_10233 = _T_6274 & _T_10232; // @[AxiLoadQueue.scala 130:72:@10541.4]
  assign _T_10235 = offsetQ_10 < 4'h9; // @[AxiLoadQueue.scala 131:33:@10542.4]
  assign _T_10238 = _T_10235 & _T_6283; // @[AxiLoadQueue.scala 131:41:@10544.4]
  assign _T_10240 = _T_10238 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10545.4]
  assign storesToCheck_10_9 = _T_2534 ? _T_10233 : _T_10240; // @[AxiLoadQueue.scala 130:10:@10546.4]
  assign _T_10246 = 4'ha <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10549.4]
  assign _T_10247 = _T_6291 & _T_10246; // @[AxiLoadQueue.scala 130:72:@10550.4]
  assign _T_10249 = offsetQ_10 < 4'ha; // @[AxiLoadQueue.scala 131:33:@10551.4]
  assign _T_10252 = _T_10249 & _T_6300; // @[AxiLoadQueue.scala 131:41:@10553.4]
  assign _T_10254 = _T_10252 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10554.4]
  assign storesToCheck_10_10 = _T_2534 ? _T_10247 : _T_10254; // @[AxiLoadQueue.scala 130:10:@10555.4]
  assign _T_10260 = 4'hb <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10558.4]
  assign _T_10261 = _T_6308 & _T_10260; // @[AxiLoadQueue.scala 130:72:@10559.4]
  assign _T_10263 = offsetQ_10 < 4'hb; // @[AxiLoadQueue.scala 131:33:@10560.4]
  assign _T_10266 = _T_10263 & _T_6317; // @[AxiLoadQueue.scala 131:41:@10562.4]
  assign _T_10268 = _T_10266 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10563.4]
  assign storesToCheck_10_11 = _T_2534 ? _T_10261 : _T_10268; // @[AxiLoadQueue.scala 130:10:@10564.4]
  assign _T_10274 = 4'hc <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10567.4]
  assign _T_10275 = _T_6325 & _T_10274; // @[AxiLoadQueue.scala 130:72:@10568.4]
  assign _T_10277 = offsetQ_10 < 4'hc; // @[AxiLoadQueue.scala 131:33:@10569.4]
  assign _T_10280 = _T_10277 & _T_6334; // @[AxiLoadQueue.scala 131:41:@10571.4]
  assign _T_10282 = _T_10280 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10572.4]
  assign storesToCheck_10_12 = _T_2534 ? _T_10275 : _T_10282; // @[AxiLoadQueue.scala 130:10:@10573.4]
  assign _T_10288 = 4'hd <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10576.4]
  assign _T_10289 = _T_6342 & _T_10288; // @[AxiLoadQueue.scala 130:72:@10577.4]
  assign _T_10291 = offsetQ_10 < 4'hd; // @[AxiLoadQueue.scala 131:33:@10578.4]
  assign _T_10294 = _T_10291 & _T_6351; // @[AxiLoadQueue.scala 131:41:@10580.4]
  assign _T_10296 = _T_10294 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10581.4]
  assign storesToCheck_10_13 = _T_2534 ? _T_10289 : _T_10296; // @[AxiLoadQueue.scala 130:10:@10582.4]
  assign _T_10302 = 4'he <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10585.4]
  assign _T_10303 = _T_6359 & _T_10302; // @[AxiLoadQueue.scala 130:72:@10586.4]
  assign _T_10305 = offsetQ_10 < 4'he; // @[AxiLoadQueue.scala 131:33:@10587.4]
  assign _T_10308 = _T_10305 & _T_6368; // @[AxiLoadQueue.scala 131:41:@10589.4]
  assign _T_10310 = _T_10308 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10590.4]
  assign storesToCheck_10_14 = _T_2534 ? _T_10303 : _T_10310; // @[AxiLoadQueue.scala 130:10:@10591.4]
  assign _T_10316 = 4'hf <= offsetQ_10; // @[AxiLoadQueue.scala 130:81:@10594.4]
  assign storesToCheck_10_15 = _T_2534 ? _T_10316 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10600.4]
  assign storesToCheck_11_0 = _T_2564 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10642.4]
  assign _T_10366 = 4'h1 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10645.4]
  assign _T_10367 = _T_6138 & _T_10366; // @[AxiLoadQueue.scala 130:72:@10646.4]
  assign _T_10369 = offsetQ_11 < 4'h1; // @[AxiLoadQueue.scala 131:33:@10647.4]
  assign _T_10372 = _T_10369 & _T_6147; // @[AxiLoadQueue.scala 131:41:@10649.4]
  assign _T_10374 = _T_10372 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10650.4]
  assign storesToCheck_11_1 = _T_2564 ? _T_10367 : _T_10374; // @[AxiLoadQueue.scala 130:10:@10651.4]
  assign _T_10380 = 4'h2 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10654.4]
  assign _T_10381 = _T_6155 & _T_10380; // @[AxiLoadQueue.scala 130:72:@10655.4]
  assign _T_10383 = offsetQ_11 < 4'h2; // @[AxiLoadQueue.scala 131:33:@10656.4]
  assign _T_10386 = _T_10383 & _T_6164; // @[AxiLoadQueue.scala 131:41:@10658.4]
  assign _T_10388 = _T_10386 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10659.4]
  assign storesToCheck_11_2 = _T_2564 ? _T_10381 : _T_10388; // @[AxiLoadQueue.scala 130:10:@10660.4]
  assign _T_10394 = 4'h3 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10663.4]
  assign _T_10395 = _T_6172 & _T_10394; // @[AxiLoadQueue.scala 130:72:@10664.4]
  assign _T_10397 = offsetQ_11 < 4'h3; // @[AxiLoadQueue.scala 131:33:@10665.4]
  assign _T_10400 = _T_10397 & _T_6181; // @[AxiLoadQueue.scala 131:41:@10667.4]
  assign _T_10402 = _T_10400 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10668.4]
  assign storesToCheck_11_3 = _T_2564 ? _T_10395 : _T_10402; // @[AxiLoadQueue.scala 130:10:@10669.4]
  assign _T_10408 = 4'h4 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10672.4]
  assign _T_10409 = _T_6189 & _T_10408; // @[AxiLoadQueue.scala 130:72:@10673.4]
  assign _T_10411 = offsetQ_11 < 4'h4; // @[AxiLoadQueue.scala 131:33:@10674.4]
  assign _T_10414 = _T_10411 & _T_6198; // @[AxiLoadQueue.scala 131:41:@10676.4]
  assign _T_10416 = _T_10414 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10677.4]
  assign storesToCheck_11_4 = _T_2564 ? _T_10409 : _T_10416; // @[AxiLoadQueue.scala 130:10:@10678.4]
  assign _T_10422 = 4'h5 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10681.4]
  assign _T_10423 = _T_6206 & _T_10422; // @[AxiLoadQueue.scala 130:72:@10682.4]
  assign _T_10425 = offsetQ_11 < 4'h5; // @[AxiLoadQueue.scala 131:33:@10683.4]
  assign _T_10428 = _T_10425 & _T_6215; // @[AxiLoadQueue.scala 131:41:@10685.4]
  assign _T_10430 = _T_10428 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10686.4]
  assign storesToCheck_11_5 = _T_2564 ? _T_10423 : _T_10430; // @[AxiLoadQueue.scala 130:10:@10687.4]
  assign _T_10436 = 4'h6 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10690.4]
  assign _T_10437 = _T_6223 & _T_10436; // @[AxiLoadQueue.scala 130:72:@10691.4]
  assign _T_10439 = offsetQ_11 < 4'h6; // @[AxiLoadQueue.scala 131:33:@10692.4]
  assign _T_10442 = _T_10439 & _T_6232; // @[AxiLoadQueue.scala 131:41:@10694.4]
  assign _T_10444 = _T_10442 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10695.4]
  assign storesToCheck_11_6 = _T_2564 ? _T_10437 : _T_10444; // @[AxiLoadQueue.scala 130:10:@10696.4]
  assign _T_10450 = 4'h7 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10699.4]
  assign _T_10451 = _T_6240 & _T_10450; // @[AxiLoadQueue.scala 130:72:@10700.4]
  assign _T_10453 = offsetQ_11 < 4'h7; // @[AxiLoadQueue.scala 131:33:@10701.4]
  assign _T_10456 = _T_10453 & _T_6249; // @[AxiLoadQueue.scala 131:41:@10703.4]
  assign _T_10458 = _T_10456 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10704.4]
  assign storesToCheck_11_7 = _T_2564 ? _T_10451 : _T_10458; // @[AxiLoadQueue.scala 130:10:@10705.4]
  assign _T_10464 = 4'h8 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10708.4]
  assign _T_10465 = _T_6257 & _T_10464; // @[AxiLoadQueue.scala 130:72:@10709.4]
  assign _T_10467 = offsetQ_11 < 4'h8; // @[AxiLoadQueue.scala 131:33:@10710.4]
  assign _T_10470 = _T_10467 & _T_6266; // @[AxiLoadQueue.scala 131:41:@10712.4]
  assign _T_10472 = _T_10470 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10713.4]
  assign storesToCheck_11_8 = _T_2564 ? _T_10465 : _T_10472; // @[AxiLoadQueue.scala 130:10:@10714.4]
  assign _T_10478 = 4'h9 <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10717.4]
  assign _T_10479 = _T_6274 & _T_10478; // @[AxiLoadQueue.scala 130:72:@10718.4]
  assign _T_10481 = offsetQ_11 < 4'h9; // @[AxiLoadQueue.scala 131:33:@10719.4]
  assign _T_10484 = _T_10481 & _T_6283; // @[AxiLoadQueue.scala 131:41:@10721.4]
  assign _T_10486 = _T_10484 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10722.4]
  assign storesToCheck_11_9 = _T_2564 ? _T_10479 : _T_10486; // @[AxiLoadQueue.scala 130:10:@10723.4]
  assign _T_10492 = 4'ha <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10726.4]
  assign _T_10493 = _T_6291 & _T_10492; // @[AxiLoadQueue.scala 130:72:@10727.4]
  assign _T_10495 = offsetQ_11 < 4'ha; // @[AxiLoadQueue.scala 131:33:@10728.4]
  assign _T_10498 = _T_10495 & _T_6300; // @[AxiLoadQueue.scala 131:41:@10730.4]
  assign _T_10500 = _T_10498 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10731.4]
  assign storesToCheck_11_10 = _T_2564 ? _T_10493 : _T_10500; // @[AxiLoadQueue.scala 130:10:@10732.4]
  assign _T_10506 = 4'hb <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10735.4]
  assign _T_10507 = _T_6308 & _T_10506; // @[AxiLoadQueue.scala 130:72:@10736.4]
  assign _T_10509 = offsetQ_11 < 4'hb; // @[AxiLoadQueue.scala 131:33:@10737.4]
  assign _T_10512 = _T_10509 & _T_6317; // @[AxiLoadQueue.scala 131:41:@10739.4]
  assign _T_10514 = _T_10512 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10740.4]
  assign storesToCheck_11_11 = _T_2564 ? _T_10507 : _T_10514; // @[AxiLoadQueue.scala 130:10:@10741.4]
  assign _T_10520 = 4'hc <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10744.4]
  assign _T_10521 = _T_6325 & _T_10520; // @[AxiLoadQueue.scala 130:72:@10745.4]
  assign _T_10523 = offsetQ_11 < 4'hc; // @[AxiLoadQueue.scala 131:33:@10746.4]
  assign _T_10526 = _T_10523 & _T_6334; // @[AxiLoadQueue.scala 131:41:@10748.4]
  assign _T_10528 = _T_10526 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10749.4]
  assign storesToCheck_11_12 = _T_2564 ? _T_10521 : _T_10528; // @[AxiLoadQueue.scala 130:10:@10750.4]
  assign _T_10534 = 4'hd <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10753.4]
  assign _T_10535 = _T_6342 & _T_10534; // @[AxiLoadQueue.scala 130:72:@10754.4]
  assign _T_10537 = offsetQ_11 < 4'hd; // @[AxiLoadQueue.scala 131:33:@10755.4]
  assign _T_10540 = _T_10537 & _T_6351; // @[AxiLoadQueue.scala 131:41:@10757.4]
  assign _T_10542 = _T_10540 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10758.4]
  assign storesToCheck_11_13 = _T_2564 ? _T_10535 : _T_10542; // @[AxiLoadQueue.scala 130:10:@10759.4]
  assign _T_10548 = 4'he <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10762.4]
  assign _T_10549 = _T_6359 & _T_10548; // @[AxiLoadQueue.scala 130:72:@10763.4]
  assign _T_10551 = offsetQ_11 < 4'he; // @[AxiLoadQueue.scala 131:33:@10764.4]
  assign _T_10554 = _T_10551 & _T_6368; // @[AxiLoadQueue.scala 131:41:@10766.4]
  assign _T_10556 = _T_10554 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10767.4]
  assign storesToCheck_11_14 = _T_2564 ? _T_10549 : _T_10556; // @[AxiLoadQueue.scala 130:10:@10768.4]
  assign _T_10562 = 4'hf <= offsetQ_11; // @[AxiLoadQueue.scala 130:81:@10771.4]
  assign storesToCheck_11_15 = _T_2564 ? _T_10562 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10777.4]
  assign storesToCheck_12_0 = _T_2594 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10819.4]
  assign _T_10612 = 4'h1 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10822.4]
  assign _T_10613 = _T_6138 & _T_10612; // @[AxiLoadQueue.scala 130:72:@10823.4]
  assign _T_10615 = offsetQ_12 < 4'h1; // @[AxiLoadQueue.scala 131:33:@10824.4]
  assign _T_10618 = _T_10615 & _T_6147; // @[AxiLoadQueue.scala 131:41:@10826.4]
  assign _T_10620 = _T_10618 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10827.4]
  assign storesToCheck_12_1 = _T_2594 ? _T_10613 : _T_10620; // @[AxiLoadQueue.scala 130:10:@10828.4]
  assign _T_10626 = 4'h2 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10831.4]
  assign _T_10627 = _T_6155 & _T_10626; // @[AxiLoadQueue.scala 130:72:@10832.4]
  assign _T_10629 = offsetQ_12 < 4'h2; // @[AxiLoadQueue.scala 131:33:@10833.4]
  assign _T_10632 = _T_10629 & _T_6164; // @[AxiLoadQueue.scala 131:41:@10835.4]
  assign _T_10634 = _T_10632 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10836.4]
  assign storesToCheck_12_2 = _T_2594 ? _T_10627 : _T_10634; // @[AxiLoadQueue.scala 130:10:@10837.4]
  assign _T_10640 = 4'h3 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10840.4]
  assign _T_10641 = _T_6172 & _T_10640; // @[AxiLoadQueue.scala 130:72:@10841.4]
  assign _T_10643 = offsetQ_12 < 4'h3; // @[AxiLoadQueue.scala 131:33:@10842.4]
  assign _T_10646 = _T_10643 & _T_6181; // @[AxiLoadQueue.scala 131:41:@10844.4]
  assign _T_10648 = _T_10646 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10845.4]
  assign storesToCheck_12_3 = _T_2594 ? _T_10641 : _T_10648; // @[AxiLoadQueue.scala 130:10:@10846.4]
  assign _T_10654 = 4'h4 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10849.4]
  assign _T_10655 = _T_6189 & _T_10654; // @[AxiLoadQueue.scala 130:72:@10850.4]
  assign _T_10657 = offsetQ_12 < 4'h4; // @[AxiLoadQueue.scala 131:33:@10851.4]
  assign _T_10660 = _T_10657 & _T_6198; // @[AxiLoadQueue.scala 131:41:@10853.4]
  assign _T_10662 = _T_10660 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10854.4]
  assign storesToCheck_12_4 = _T_2594 ? _T_10655 : _T_10662; // @[AxiLoadQueue.scala 130:10:@10855.4]
  assign _T_10668 = 4'h5 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10858.4]
  assign _T_10669 = _T_6206 & _T_10668; // @[AxiLoadQueue.scala 130:72:@10859.4]
  assign _T_10671 = offsetQ_12 < 4'h5; // @[AxiLoadQueue.scala 131:33:@10860.4]
  assign _T_10674 = _T_10671 & _T_6215; // @[AxiLoadQueue.scala 131:41:@10862.4]
  assign _T_10676 = _T_10674 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10863.4]
  assign storesToCheck_12_5 = _T_2594 ? _T_10669 : _T_10676; // @[AxiLoadQueue.scala 130:10:@10864.4]
  assign _T_10682 = 4'h6 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10867.4]
  assign _T_10683 = _T_6223 & _T_10682; // @[AxiLoadQueue.scala 130:72:@10868.4]
  assign _T_10685 = offsetQ_12 < 4'h6; // @[AxiLoadQueue.scala 131:33:@10869.4]
  assign _T_10688 = _T_10685 & _T_6232; // @[AxiLoadQueue.scala 131:41:@10871.4]
  assign _T_10690 = _T_10688 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10872.4]
  assign storesToCheck_12_6 = _T_2594 ? _T_10683 : _T_10690; // @[AxiLoadQueue.scala 130:10:@10873.4]
  assign _T_10696 = 4'h7 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10876.4]
  assign _T_10697 = _T_6240 & _T_10696; // @[AxiLoadQueue.scala 130:72:@10877.4]
  assign _T_10699 = offsetQ_12 < 4'h7; // @[AxiLoadQueue.scala 131:33:@10878.4]
  assign _T_10702 = _T_10699 & _T_6249; // @[AxiLoadQueue.scala 131:41:@10880.4]
  assign _T_10704 = _T_10702 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10881.4]
  assign storesToCheck_12_7 = _T_2594 ? _T_10697 : _T_10704; // @[AxiLoadQueue.scala 130:10:@10882.4]
  assign _T_10710 = 4'h8 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10885.4]
  assign _T_10711 = _T_6257 & _T_10710; // @[AxiLoadQueue.scala 130:72:@10886.4]
  assign _T_10713 = offsetQ_12 < 4'h8; // @[AxiLoadQueue.scala 131:33:@10887.4]
  assign _T_10716 = _T_10713 & _T_6266; // @[AxiLoadQueue.scala 131:41:@10889.4]
  assign _T_10718 = _T_10716 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10890.4]
  assign storesToCheck_12_8 = _T_2594 ? _T_10711 : _T_10718; // @[AxiLoadQueue.scala 130:10:@10891.4]
  assign _T_10724 = 4'h9 <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10894.4]
  assign _T_10725 = _T_6274 & _T_10724; // @[AxiLoadQueue.scala 130:72:@10895.4]
  assign _T_10727 = offsetQ_12 < 4'h9; // @[AxiLoadQueue.scala 131:33:@10896.4]
  assign _T_10730 = _T_10727 & _T_6283; // @[AxiLoadQueue.scala 131:41:@10898.4]
  assign _T_10732 = _T_10730 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10899.4]
  assign storesToCheck_12_9 = _T_2594 ? _T_10725 : _T_10732; // @[AxiLoadQueue.scala 130:10:@10900.4]
  assign _T_10738 = 4'ha <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10903.4]
  assign _T_10739 = _T_6291 & _T_10738; // @[AxiLoadQueue.scala 130:72:@10904.4]
  assign _T_10741 = offsetQ_12 < 4'ha; // @[AxiLoadQueue.scala 131:33:@10905.4]
  assign _T_10744 = _T_10741 & _T_6300; // @[AxiLoadQueue.scala 131:41:@10907.4]
  assign _T_10746 = _T_10744 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10908.4]
  assign storesToCheck_12_10 = _T_2594 ? _T_10739 : _T_10746; // @[AxiLoadQueue.scala 130:10:@10909.4]
  assign _T_10752 = 4'hb <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10912.4]
  assign _T_10753 = _T_6308 & _T_10752; // @[AxiLoadQueue.scala 130:72:@10913.4]
  assign _T_10755 = offsetQ_12 < 4'hb; // @[AxiLoadQueue.scala 131:33:@10914.4]
  assign _T_10758 = _T_10755 & _T_6317; // @[AxiLoadQueue.scala 131:41:@10916.4]
  assign _T_10760 = _T_10758 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10917.4]
  assign storesToCheck_12_11 = _T_2594 ? _T_10753 : _T_10760; // @[AxiLoadQueue.scala 130:10:@10918.4]
  assign _T_10766 = 4'hc <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10921.4]
  assign _T_10767 = _T_6325 & _T_10766; // @[AxiLoadQueue.scala 130:72:@10922.4]
  assign _T_10769 = offsetQ_12 < 4'hc; // @[AxiLoadQueue.scala 131:33:@10923.4]
  assign _T_10772 = _T_10769 & _T_6334; // @[AxiLoadQueue.scala 131:41:@10925.4]
  assign _T_10774 = _T_10772 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10926.4]
  assign storesToCheck_12_12 = _T_2594 ? _T_10767 : _T_10774; // @[AxiLoadQueue.scala 130:10:@10927.4]
  assign _T_10780 = 4'hd <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10930.4]
  assign _T_10781 = _T_6342 & _T_10780; // @[AxiLoadQueue.scala 130:72:@10931.4]
  assign _T_10783 = offsetQ_12 < 4'hd; // @[AxiLoadQueue.scala 131:33:@10932.4]
  assign _T_10786 = _T_10783 & _T_6351; // @[AxiLoadQueue.scala 131:41:@10934.4]
  assign _T_10788 = _T_10786 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10935.4]
  assign storesToCheck_12_13 = _T_2594 ? _T_10781 : _T_10788; // @[AxiLoadQueue.scala 130:10:@10936.4]
  assign _T_10794 = 4'he <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10939.4]
  assign _T_10795 = _T_6359 & _T_10794; // @[AxiLoadQueue.scala 130:72:@10940.4]
  assign _T_10797 = offsetQ_12 < 4'he; // @[AxiLoadQueue.scala 131:33:@10941.4]
  assign _T_10800 = _T_10797 & _T_6368; // @[AxiLoadQueue.scala 131:41:@10943.4]
  assign _T_10802 = _T_10800 == 1'h0; // @[AxiLoadQueue.scala 131:9:@10944.4]
  assign storesToCheck_12_14 = _T_2594 ? _T_10795 : _T_10802; // @[AxiLoadQueue.scala 130:10:@10945.4]
  assign _T_10808 = 4'hf <= offsetQ_12; // @[AxiLoadQueue.scala 130:81:@10948.4]
  assign storesToCheck_12_15 = _T_2594 ? _T_10808 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10954.4]
  assign storesToCheck_13_0 = _T_2624 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@10996.4]
  assign _T_10858 = 4'h1 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@10999.4]
  assign _T_10859 = _T_6138 & _T_10858; // @[AxiLoadQueue.scala 130:72:@11000.4]
  assign _T_10861 = offsetQ_13 < 4'h1; // @[AxiLoadQueue.scala 131:33:@11001.4]
  assign _T_10864 = _T_10861 & _T_6147; // @[AxiLoadQueue.scala 131:41:@11003.4]
  assign _T_10866 = _T_10864 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11004.4]
  assign storesToCheck_13_1 = _T_2624 ? _T_10859 : _T_10866; // @[AxiLoadQueue.scala 130:10:@11005.4]
  assign _T_10872 = 4'h2 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11008.4]
  assign _T_10873 = _T_6155 & _T_10872; // @[AxiLoadQueue.scala 130:72:@11009.4]
  assign _T_10875 = offsetQ_13 < 4'h2; // @[AxiLoadQueue.scala 131:33:@11010.4]
  assign _T_10878 = _T_10875 & _T_6164; // @[AxiLoadQueue.scala 131:41:@11012.4]
  assign _T_10880 = _T_10878 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11013.4]
  assign storesToCheck_13_2 = _T_2624 ? _T_10873 : _T_10880; // @[AxiLoadQueue.scala 130:10:@11014.4]
  assign _T_10886 = 4'h3 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11017.4]
  assign _T_10887 = _T_6172 & _T_10886; // @[AxiLoadQueue.scala 130:72:@11018.4]
  assign _T_10889 = offsetQ_13 < 4'h3; // @[AxiLoadQueue.scala 131:33:@11019.4]
  assign _T_10892 = _T_10889 & _T_6181; // @[AxiLoadQueue.scala 131:41:@11021.4]
  assign _T_10894 = _T_10892 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11022.4]
  assign storesToCheck_13_3 = _T_2624 ? _T_10887 : _T_10894; // @[AxiLoadQueue.scala 130:10:@11023.4]
  assign _T_10900 = 4'h4 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11026.4]
  assign _T_10901 = _T_6189 & _T_10900; // @[AxiLoadQueue.scala 130:72:@11027.4]
  assign _T_10903 = offsetQ_13 < 4'h4; // @[AxiLoadQueue.scala 131:33:@11028.4]
  assign _T_10906 = _T_10903 & _T_6198; // @[AxiLoadQueue.scala 131:41:@11030.4]
  assign _T_10908 = _T_10906 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11031.4]
  assign storesToCheck_13_4 = _T_2624 ? _T_10901 : _T_10908; // @[AxiLoadQueue.scala 130:10:@11032.4]
  assign _T_10914 = 4'h5 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11035.4]
  assign _T_10915 = _T_6206 & _T_10914; // @[AxiLoadQueue.scala 130:72:@11036.4]
  assign _T_10917 = offsetQ_13 < 4'h5; // @[AxiLoadQueue.scala 131:33:@11037.4]
  assign _T_10920 = _T_10917 & _T_6215; // @[AxiLoadQueue.scala 131:41:@11039.4]
  assign _T_10922 = _T_10920 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11040.4]
  assign storesToCheck_13_5 = _T_2624 ? _T_10915 : _T_10922; // @[AxiLoadQueue.scala 130:10:@11041.4]
  assign _T_10928 = 4'h6 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11044.4]
  assign _T_10929 = _T_6223 & _T_10928; // @[AxiLoadQueue.scala 130:72:@11045.4]
  assign _T_10931 = offsetQ_13 < 4'h6; // @[AxiLoadQueue.scala 131:33:@11046.4]
  assign _T_10934 = _T_10931 & _T_6232; // @[AxiLoadQueue.scala 131:41:@11048.4]
  assign _T_10936 = _T_10934 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11049.4]
  assign storesToCheck_13_6 = _T_2624 ? _T_10929 : _T_10936; // @[AxiLoadQueue.scala 130:10:@11050.4]
  assign _T_10942 = 4'h7 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11053.4]
  assign _T_10943 = _T_6240 & _T_10942; // @[AxiLoadQueue.scala 130:72:@11054.4]
  assign _T_10945 = offsetQ_13 < 4'h7; // @[AxiLoadQueue.scala 131:33:@11055.4]
  assign _T_10948 = _T_10945 & _T_6249; // @[AxiLoadQueue.scala 131:41:@11057.4]
  assign _T_10950 = _T_10948 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11058.4]
  assign storesToCheck_13_7 = _T_2624 ? _T_10943 : _T_10950; // @[AxiLoadQueue.scala 130:10:@11059.4]
  assign _T_10956 = 4'h8 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11062.4]
  assign _T_10957 = _T_6257 & _T_10956; // @[AxiLoadQueue.scala 130:72:@11063.4]
  assign _T_10959 = offsetQ_13 < 4'h8; // @[AxiLoadQueue.scala 131:33:@11064.4]
  assign _T_10962 = _T_10959 & _T_6266; // @[AxiLoadQueue.scala 131:41:@11066.4]
  assign _T_10964 = _T_10962 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11067.4]
  assign storesToCheck_13_8 = _T_2624 ? _T_10957 : _T_10964; // @[AxiLoadQueue.scala 130:10:@11068.4]
  assign _T_10970 = 4'h9 <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11071.4]
  assign _T_10971 = _T_6274 & _T_10970; // @[AxiLoadQueue.scala 130:72:@11072.4]
  assign _T_10973 = offsetQ_13 < 4'h9; // @[AxiLoadQueue.scala 131:33:@11073.4]
  assign _T_10976 = _T_10973 & _T_6283; // @[AxiLoadQueue.scala 131:41:@11075.4]
  assign _T_10978 = _T_10976 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11076.4]
  assign storesToCheck_13_9 = _T_2624 ? _T_10971 : _T_10978; // @[AxiLoadQueue.scala 130:10:@11077.4]
  assign _T_10984 = 4'ha <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11080.4]
  assign _T_10985 = _T_6291 & _T_10984; // @[AxiLoadQueue.scala 130:72:@11081.4]
  assign _T_10987 = offsetQ_13 < 4'ha; // @[AxiLoadQueue.scala 131:33:@11082.4]
  assign _T_10990 = _T_10987 & _T_6300; // @[AxiLoadQueue.scala 131:41:@11084.4]
  assign _T_10992 = _T_10990 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11085.4]
  assign storesToCheck_13_10 = _T_2624 ? _T_10985 : _T_10992; // @[AxiLoadQueue.scala 130:10:@11086.4]
  assign _T_10998 = 4'hb <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11089.4]
  assign _T_10999 = _T_6308 & _T_10998; // @[AxiLoadQueue.scala 130:72:@11090.4]
  assign _T_11001 = offsetQ_13 < 4'hb; // @[AxiLoadQueue.scala 131:33:@11091.4]
  assign _T_11004 = _T_11001 & _T_6317; // @[AxiLoadQueue.scala 131:41:@11093.4]
  assign _T_11006 = _T_11004 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11094.4]
  assign storesToCheck_13_11 = _T_2624 ? _T_10999 : _T_11006; // @[AxiLoadQueue.scala 130:10:@11095.4]
  assign _T_11012 = 4'hc <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11098.4]
  assign _T_11013 = _T_6325 & _T_11012; // @[AxiLoadQueue.scala 130:72:@11099.4]
  assign _T_11015 = offsetQ_13 < 4'hc; // @[AxiLoadQueue.scala 131:33:@11100.4]
  assign _T_11018 = _T_11015 & _T_6334; // @[AxiLoadQueue.scala 131:41:@11102.4]
  assign _T_11020 = _T_11018 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11103.4]
  assign storesToCheck_13_12 = _T_2624 ? _T_11013 : _T_11020; // @[AxiLoadQueue.scala 130:10:@11104.4]
  assign _T_11026 = 4'hd <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11107.4]
  assign _T_11027 = _T_6342 & _T_11026; // @[AxiLoadQueue.scala 130:72:@11108.4]
  assign _T_11029 = offsetQ_13 < 4'hd; // @[AxiLoadQueue.scala 131:33:@11109.4]
  assign _T_11032 = _T_11029 & _T_6351; // @[AxiLoadQueue.scala 131:41:@11111.4]
  assign _T_11034 = _T_11032 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11112.4]
  assign storesToCheck_13_13 = _T_2624 ? _T_11027 : _T_11034; // @[AxiLoadQueue.scala 130:10:@11113.4]
  assign _T_11040 = 4'he <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11116.4]
  assign _T_11041 = _T_6359 & _T_11040; // @[AxiLoadQueue.scala 130:72:@11117.4]
  assign _T_11043 = offsetQ_13 < 4'he; // @[AxiLoadQueue.scala 131:33:@11118.4]
  assign _T_11046 = _T_11043 & _T_6368; // @[AxiLoadQueue.scala 131:41:@11120.4]
  assign _T_11048 = _T_11046 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11121.4]
  assign storesToCheck_13_14 = _T_2624 ? _T_11041 : _T_11048; // @[AxiLoadQueue.scala 130:10:@11122.4]
  assign _T_11054 = 4'hf <= offsetQ_13; // @[AxiLoadQueue.scala 130:81:@11125.4]
  assign storesToCheck_13_15 = _T_2624 ? _T_11054 : 1'h1; // @[AxiLoadQueue.scala 130:10:@11131.4]
  assign storesToCheck_14_0 = _T_2654 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@11173.4]
  assign _T_11104 = 4'h1 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11176.4]
  assign _T_11105 = _T_6138 & _T_11104; // @[AxiLoadQueue.scala 130:72:@11177.4]
  assign _T_11107 = offsetQ_14 < 4'h1; // @[AxiLoadQueue.scala 131:33:@11178.4]
  assign _T_11110 = _T_11107 & _T_6147; // @[AxiLoadQueue.scala 131:41:@11180.4]
  assign _T_11112 = _T_11110 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11181.4]
  assign storesToCheck_14_1 = _T_2654 ? _T_11105 : _T_11112; // @[AxiLoadQueue.scala 130:10:@11182.4]
  assign _T_11118 = 4'h2 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11185.4]
  assign _T_11119 = _T_6155 & _T_11118; // @[AxiLoadQueue.scala 130:72:@11186.4]
  assign _T_11121 = offsetQ_14 < 4'h2; // @[AxiLoadQueue.scala 131:33:@11187.4]
  assign _T_11124 = _T_11121 & _T_6164; // @[AxiLoadQueue.scala 131:41:@11189.4]
  assign _T_11126 = _T_11124 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11190.4]
  assign storesToCheck_14_2 = _T_2654 ? _T_11119 : _T_11126; // @[AxiLoadQueue.scala 130:10:@11191.4]
  assign _T_11132 = 4'h3 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11194.4]
  assign _T_11133 = _T_6172 & _T_11132; // @[AxiLoadQueue.scala 130:72:@11195.4]
  assign _T_11135 = offsetQ_14 < 4'h3; // @[AxiLoadQueue.scala 131:33:@11196.4]
  assign _T_11138 = _T_11135 & _T_6181; // @[AxiLoadQueue.scala 131:41:@11198.4]
  assign _T_11140 = _T_11138 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11199.4]
  assign storesToCheck_14_3 = _T_2654 ? _T_11133 : _T_11140; // @[AxiLoadQueue.scala 130:10:@11200.4]
  assign _T_11146 = 4'h4 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11203.4]
  assign _T_11147 = _T_6189 & _T_11146; // @[AxiLoadQueue.scala 130:72:@11204.4]
  assign _T_11149 = offsetQ_14 < 4'h4; // @[AxiLoadQueue.scala 131:33:@11205.4]
  assign _T_11152 = _T_11149 & _T_6198; // @[AxiLoadQueue.scala 131:41:@11207.4]
  assign _T_11154 = _T_11152 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11208.4]
  assign storesToCheck_14_4 = _T_2654 ? _T_11147 : _T_11154; // @[AxiLoadQueue.scala 130:10:@11209.4]
  assign _T_11160 = 4'h5 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11212.4]
  assign _T_11161 = _T_6206 & _T_11160; // @[AxiLoadQueue.scala 130:72:@11213.4]
  assign _T_11163 = offsetQ_14 < 4'h5; // @[AxiLoadQueue.scala 131:33:@11214.4]
  assign _T_11166 = _T_11163 & _T_6215; // @[AxiLoadQueue.scala 131:41:@11216.4]
  assign _T_11168 = _T_11166 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11217.4]
  assign storesToCheck_14_5 = _T_2654 ? _T_11161 : _T_11168; // @[AxiLoadQueue.scala 130:10:@11218.4]
  assign _T_11174 = 4'h6 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11221.4]
  assign _T_11175 = _T_6223 & _T_11174; // @[AxiLoadQueue.scala 130:72:@11222.4]
  assign _T_11177 = offsetQ_14 < 4'h6; // @[AxiLoadQueue.scala 131:33:@11223.4]
  assign _T_11180 = _T_11177 & _T_6232; // @[AxiLoadQueue.scala 131:41:@11225.4]
  assign _T_11182 = _T_11180 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11226.4]
  assign storesToCheck_14_6 = _T_2654 ? _T_11175 : _T_11182; // @[AxiLoadQueue.scala 130:10:@11227.4]
  assign _T_11188 = 4'h7 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11230.4]
  assign _T_11189 = _T_6240 & _T_11188; // @[AxiLoadQueue.scala 130:72:@11231.4]
  assign _T_11191 = offsetQ_14 < 4'h7; // @[AxiLoadQueue.scala 131:33:@11232.4]
  assign _T_11194 = _T_11191 & _T_6249; // @[AxiLoadQueue.scala 131:41:@11234.4]
  assign _T_11196 = _T_11194 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11235.4]
  assign storesToCheck_14_7 = _T_2654 ? _T_11189 : _T_11196; // @[AxiLoadQueue.scala 130:10:@11236.4]
  assign _T_11202 = 4'h8 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11239.4]
  assign _T_11203 = _T_6257 & _T_11202; // @[AxiLoadQueue.scala 130:72:@11240.4]
  assign _T_11205 = offsetQ_14 < 4'h8; // @[AxiLoadQueue.scala 131:33:@11241.4]
  assign _T_11208 = _T_11205 & _T_6266; // @[AxiLoadQueue.scala 131:41:@11243.4]
  assign _T_11210 = _T_11208 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11244.4]
  assign storesToCheck_14_8 = _T_2654 ? _T_11203 : _T_11210; // @[AxiLoadQueue.scala 130:10:@11245.4]
  assign _T_11216 = 4'h9 <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11248.4]
  assign _T_11217 = _T_6274 & _T_11216; // @[AxiLoadQueue.scala 130:72:@11249.4]
  assign _T_11219 = offsetQ_14 < 4'h9; // @[AxiLoadQueue.scala 131:33:@11250.4]
  assign _T_11222 = _T_11219 & _T_6283; // @[AxiLoadQueue.scala 131:41:@11252.4]
  assign _T_11224 = _T_11222 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11253.4]
  assign storesToCheck_14_9 = _T_2654 ? _T_11217 : _T_11224; // @[AxiLoadQueue.scala 130:10:@11254.4]
  assign _T_11230 = 4'ha <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11257.4]
  assign _T_11231 = _T_6291 & _T_11230; // @[AxiLoadQueue.scala 130:72:@11258.4]
  assign _T_11233 = offsetQ_14 < 4'ha; // @[AxiLoadQueue.scala 131:33:@11259.4]
  assign _T_11236 = _T_11233 & _T_6300; // @[AxiLoadQueue.scala 131:41:@11261.4]
  assign _T_11238 = _T_11236 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11262.4]
  assign storesToCheck_14_10 = _T_2654 ? _T_11231 : _T_11238; // @[AxiLoadQueue.scala 130:10:@11263.4]
  assign _T_11244 = 4'hb <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11266.4]
  assign _T_11245 = _T_6308 & _T_11244; // @[AxiLoadQueue.scala 130:72:@11267.4]
  assign _T_11247 = offsetQ_14 < 4'hb; // @[AxiLoadQueue.scala 131:33:@11268.4]
  assign _T_11250 = _T_11247 & _T_6317; // @[AxiLoadQueue.scala 131:41:@11270.4]
  assign _T_11252 = _T_11250 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11271.4]
  assign storesToCheck_14_11 = _T_2654 ? _T_11245 : _T_11252; // @[AxiLoadQueue.scala 130:10:@11272.4]
  assign _T_11258 = 4'hc <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11275.4]
  assign _T_11259 = _T_6325 & _T_11258; // @[AxiLoadQueue.scala 130:72:@11276.4]
  assign _T_11261 = offsetQ_14 < 4'hc; // @[AxiLoadQueue.scala 131:33:@11277.4]
  assign _T_11264 = _T_11261 & _T_6334; // @[AxiLoadQueue.scala 131:41:@11279.4]
  assign _T_11266 = _T_11264 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11280.4]
  assign storesToCheck_14_12 = _T_2654 ? _T_11259 : _T_11266; // @[AxiLoadQueue.scala 130:10:@11281.4]
  assign _T_11272 = 4'hd <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11284.4]
  assign _T_11273 = _T_6342 & _T_11272; // @[AxiLoadQueue.scala 130:72:@11285.4]
  assign _T_11275 = offsetQ_14 < 4'hd; // @[AxiLoadQueue.scala 131:33:@11286.4]
  assign _T_11278 = _T_11275 & _T_6351; // @[AxiLoadQueue.scala 131:41:@11288.4]
  assign _T_11280 = _T_11278 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11289.4]
  assign storesToCheck_14_13 = _T_2654 ? _T_11273 : _T_11280; // @[AxiLoadQueue.scala 130:10:@11290.4]
  assign _T_11286 = 4'he <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11293.4]
  assign _T_11287 = _T_6359 & _T_11286; // @[AxiLoadQueue.scala 130:72:@11294.4]
  assign _T_11289 = offsetQ_14 < 4'he; // @[AxiLoadQueue.scala 131:33:@11295.4]
  assign _T_11292 = _T_11289 & _T_6368; // @[AxiLoadQueue.scala 131:41:@11297.4]
  assign _T_11294 = _T_11292 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11298.4]
  assign storesToCheck_14_14 = _T_2654 ? _T_11287 : _T_11294; // @[AxiLoadQueue.scala 130:10:@11299.4]
  assign _T_11300 = 4'hf <= offsetQ_14; // @[AxiLoadQueue.scala 130:81:@11302.4]
  assign storesToCheck_14_15 = _T_2654 ? _T_11300 : 1'h1; // @[AxiLoadQueue.scala 130:10:@11308.4]
  assign storesToCheck_15_0 = _T_2684 ? _T_6121 : 1'h1; // @[AxiLoadQueue.scala 130:10:@11350.4]
  assign _T_11350 = 4'h1 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11353.4]
  assign _T_11351 = _T_6138 & _T_11350; // @[AxiLoadQueue.scala 130:72:@11354.4]
  assign _T_11353 = offsetQ_15 < 4'h1; // @[AxiLoadQueue.scala 131:33:@11355.4]
  assign _T_11356 = _T_11353 & _T_6147; // @[AxiLoadQueue.scala 131:41:@11357.4]
  assign _T_11358 = _T_11356 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11358.4]
  assign storesToCheck_15_1 = _T_2684 ? _T_11351 : _T_11358; // @[AxiLoadQueue.scala 130:10:@11359.4]
  assign _T_11364 = 4'h2 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11362.4]
  assign _T_11365 = _T_6155 & _T_11364; // @[AxiLoadQueue.scala 130:72:@11363.4]
  assign _T_11367 = offsetQ_15 < 4'h2; // @[AxiLoadQueue.scala 131:33:@11364.4]
  assign _T_11370 = _T_11367 & _T_6164; // @[AxiLoadQueue.scala 131:41:@11366.4]
  assign _T_11372 = _T_11370 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11367.4]
  assign storesToCheck_15_2 = _T_2684 ? _T_11365 : _T_11372; // @[AxiLoadQueue.scala 130:10:@11368.4]
  assign _T_11378 = 4'h3 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11371.4]
  assign _T_11379 = _T_6172 & _T_11378; // @[AxiLoadQueue.scala 130:72:@11372.4]
  assign _T_11381 = offsetQ_15 < 4'h3; // @[AxiLoadQueue.scala 131:33:@11373.4]
  assign _T_11384 = _T_11381 & _T_6181; // @[AxiLoadQueue.scala 131:41:@11375.4]
  assign _T_11386 = _T_11384 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11376.4]
  assign storesToCheck_15_3 = _T_2684 ? _T_11379 : _T_11386; // @[AxiLoadQueue.scala 130:10:@11377.4]
  assign _T_11392 = 4'h4 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11380.4]
  assign _T_11393 = _T_6189 & _T_11392; // @[AxiLoadQueue.scala 130:72:@11381.4]
  assign _T_11395 = offsetQ_15 < 4'h4; // @[AxiLoadQueue.scala 131:33:@11382.4]
  assign _T_11398 = _T_11395 & _T_6198; // @[AxiLoadQueue.scala 131:41:@11384.4]
  assign _T_11400 = _T_11398 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11385.4]
  assign storesToCheck_15_4 = _T_2684 ? _T_11393 : _T_11400; // @[AxiLoadQueue.scala 130:10:@11386.4]
  assign _T_11406 = 4'h5 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11389.4]
  assign _T_11407 = _T_6206 & _T_11406; // @[AxiLoadQueue.scala 130:72:@11390.4]
  assign _T_11409 = offsetQ_15 < 4'h5; // @[AxiLoadQueue.scala 131:33:@11391.4]
  assign _T_11412 = _T_11409 & _T_6215; // @[AxiLoadQueue.scala 131:41:@11393.4]
  assign _T_11414 = _T_11412 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11394.4]
  assign storesToCheck_15_5 = _T_2684 ? _T_11407 : _T_11414; // @[AxiLoadQueue.scala 130:10:@11395.4]
  assign _T_11420 = 4'h6 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11398.4]
  assign _T_11421 = _T_6223 & _T_11420; // @[AxiLoadQueue.scala 130:72:@11399.4]
  assign _T_11423 = offsetQ_15 < 4'h6; // @[AxiLoadQueue.scala 131:33:@11400.4]
  assign _T_11426 = _T_11423 & _T_6232; // @[AxiLoadQueue.scala 131:41:@11402.4]
  assign _T_11428 = _T_11426 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11403.4]
  assign storesToCheck_15_6 = _T_2684 ? _T_11421 : _T_11428; // @[AxiLoadQueue.scala 130:10:@11404.4]
  assign _T_11434 = 4'h7 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11407.4]
  assign _T_11435 = _T_6240 & _T_11434; // @[AxiLoadQueue.scala 130:72:@11408.4]
  assign _T_11437 = offsetQ_15 < 4'h7; // @[AxiLoadQueue.scala 131:33:@11409.4]
  assign _T_11440 = _T_11437 & _T_6249; // @[AxiLoadQueue.scala 131:41:@11411.4]
  assign _T_11442 = _T_11440 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11412.4]
  assign storesToCheck_15_7 = _T_2684 ? _T_11435 : _T_11442; // @[AxiLoadQueue.scala 130:10:@11413.4]
  assign _T_11448 = 4'h8 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11416.4]
  assign _T_11449 = _T_6257 & _T_11448; // @[AxiLoadQueue.scala 130:72:@11417.4]
  assign _T_11451 = offsetQ_15 < 4'h8; // @[AxiLoadQueue.scala 131:33:@11418.4]
  assign _T_11454 = _T_11451 & _T_6266; // @[AxiLoadQueue.scala 131:41:@11420.4]
  assign _T_11456 = _T_11454 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11421.4]
  assign storesToCheck_15_8 = _T_2684 ? _T_11449 : _T_11456; // @[AxiLoadQueue.scala 130:10:@11422.4]
  assign _T_11462 = 4'h9 <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11425.4]
  assign _T_11463 = _T_6274 & _T_11462; // @[AxiLoadQueue.scala 130:72:@11426.4]
  assign _T_11465 = offsetQ_15 < 4'h9; // @[AxiLoadQueue.scala 131:33:@11427.4]
  assign _T_11468 = _T_11465 & _T_6283; // @[AxiLoadQueue.scala 131:41:@11429.4]
  assign _T_11470 = _T_11468 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11430.4]
  assign storesToCheck_15_9 = _T_2684 ? _T_11463 : _T_11470; // @[AxiLoadQueue.scala 130:10:@11431.4]
  assign _T_11476 = 4'ha <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11434.4]
  assign _T_11477 = _T_6291 & _T_11476; // @[AxiLoadQueue.scala 130:72:@11435.4]
  assign _T_11479 = offsetQ_15 < 4'ha; // @[AxiLoadQueue.scala 131:33:@11436.4]
  assign _T_11482 = _T_11479 & _T_6300; // @[AxiLoadQueue.scala 131:41:@11438.4]
  assign _T_11484 = _T_11482 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11439.4]
  assign storesToCheck_15_10 = _T_2684 ? _T_11477 : _T_11484; // @[AxiLoadQueue.scala 130:10:@11440.4]
  assign _T_11490 = 4'hb <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11443.4]
  assign _T_11491 = _T_6308 & _T_11490; // @[AxiLoadQueue.scala 130:72:@11444.4]
  assign _T_11493 = offsetQ_15 < 4'hb; // @[AxiLoadQueue.scala 131:33:@11445.4]
  assign _T_11496 = _T_11493 & _T_6317; // @[AxiLoadQueue.scala 131:41:@11447.4]
  assign _T_11498 = _T_11496 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11448.4]
  assign storesToCheck_15_11 = _T_2684 ? _T_11491 : _T_11498; // @[AxiLoadQueue.scala 130:10:@11449.4]
  assign _T_11504 = 4'hc <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11452.4]
  assign _T_11505 = _T_6325 & _T_11504; // @[AxiLoadQueue.scala 130:72:@11453.4]
  assign _T_11507 = offsetQ_15 < 4'hc; // @[AxiLoadQueue.scala 131:33:@11454.4]
  assign _T_11510 = _T_11507 & _T_6334; // @[AxiLoadQueue.scala 131:41:@11456.4]
  assign _T_11512 = _T_11510 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11457.4]
  assign storesToCheck_15_12 = _T_2684 ? _T_11505 : _T_11512; // @[AxiLoadQueue.scala 130:10:@11458.4]
  assign _T_11518 = 4'hd <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11461.4]
  assign _T_11519 = _T_6342 & _T_11518; // @[AxiLoadQueue.scala 130:72:@11462.4]
  assign _T_11521 = offsetQ_15 < 4'hd; // @[AxiLoadQueue.scala 131:33:@11463.4]
  assign _T_11524 = _T_11521 & _T_6351; // @[AxiLoadQueue.scala 131:41:@11465.4]
  assign _T_11526 = _T_11524 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11466.4]
  assign storesToCheck_15_13 = _T_2684 ? _T_11519 : _T_11526; // @[AxiLoadQueue.scala 130:10:@11467.4]
  assign _T_11532 = 4'he <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11470.4]
  assign _T_11533 = _T_6359 & _T_11532; // @[AxiLoadQueue.scala 130:72:@11471.4]
  assign _T_11535 = offsetQ_15 < 4'he; // @[AxiLoadQueue.scala 131:33:@11472.4]
  assign _T_11538 = _T_11535 & _T_6368; // @[AxiLoadQueue.scala 131:41:@11474.4]
  assign _T_11540 = _T_11538 == 1'h0; // @[AxiLoadQueue.scala 131:9:@11475.4]
  assign storesToCheck_15_14 = _T_2684 ? _T_11533 : _T_11540; // @[AxiLoadQueue.scala 130:10:@11476.4]
  assign _T_11546 = 4'hf <= offsetQ_15; // @[AxiLoadQueue.scala 130:81:@11479.4]
  assign storesToCheck_15_15 = _T_2684 ? _T_11546 : 1'h1; // @[AxiLoadQueue.scala 130:10:@11485.4]
  assign _T_12808 = storesToCheck_0_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11520.4]
  assign entriesToCheck_0_0 = _T_12808 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11521.4]
  assign _T_12810 = storesToCheck_0_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11522.4]
  assign entriesToCheck_0_1 = _T_12810 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11523.4]
  assign _T_12812 = storesToCheck_0_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11524.4]
  assign entriesToCheck_0_2 = _T_12812 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11525.4]
  assign _T_12814 = storesToCheck_0_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11526.4]
  assign entriesToCheck_0_3 = _T_12814 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11527.4]
  assign _T_12816 = storesToCheck_0_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11528.4]
  assign entriesToCheck_0_4 = _T_12816 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11529.4]
  assign _T_12818 = storesToCheck_0_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11530.4]
  assign entriesToCheck_0_5 = _T_12818 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11531.4]
  assign _T_12820 = storesToCheck_0_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11532.4]
  assign entriesToCheck_0_6 = _T_12820 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11533.4]
  assign _T_12822 = storesToCheck_0_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11534.4]
  assign entriesToCheck_0_7 = _T_12822 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11535.4]
  assign _T_12824 = storesToCheck_0_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11536.4]
  assign entriesToCheck_0_8 = _T_12824 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11537.4]
  assign _T_12826 = storesToCheck_0_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11538.4]
  assign entriesToCheck_0_9 = _T_12826 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11539.4]
  assign _T_12828 = storesToCheck_0_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11540.4]
  assign entriesToCheck_0_10 = _T_12828 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11541.4]
  assign _T_12830 = storesToCheck_0_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11542.4]
  assign entriesToCheck_0_11 = _T_12830 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11543.4]
  assign _T_12832 = storesToCheck_0_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11544.4]
  assign entriesToCheck_0_12 = _T_12832 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11545.4]
  assign _T_12834 = storesToCheck_0_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11546.4]
  assign entriesToCheck_0_13 = _T_12834 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11547.4]
  assign _T_12836 = storesToCheck_0_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11548.4]
  assign entriesToCheck_0_14 = _T_12836 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11549.4]
  assign _T_12838 = storesToCheck_0_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11550.4]
  assign entriesToCheck_0_15 = _T_12838 & checkBits_0; // @[AxiLoadQueue.scala 140:26:@11551.4]
  assign _T_12840 = storesToCheck_1_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11568.4]
  assign entriesToCheck_1_0 = _T_12840 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11569.4]
  assign _T_12842 = storesToCheck_1_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11570.4]
  assign entriesToCheck_1_1 = _T_12842 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11571.4]
  assign _T_12844 = storesToCheck_1_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11572.4]
  assign entriesToCheck_1_2 = _T_12844 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11573.4]
  assign _T_12846 = storesToCheck_1_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11574.4]
  assign entriesToCheck_1_3 = _T_12846 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11575.4]
  assign _T_12848 = storesToCheck_1_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11576.4]
  assign entriesToCheck_1_4 = _T_12848 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11577.4]
  assign _T_12850 = storesToCheck_1_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11578.4]
  assign entriesToCheck_1_5 = _T_12850 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11579.4]
  assign _T_12852 = storesToCheck_1_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11580.4]
  assign entriesToCheck_1_6 = _T_12852 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11581.4]
  assign _T_12854 = storesToCheck_1_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11582.4]
  assign entriesToCheck_1_7 = _T_12854 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11583.4]
  assign _T_12856 = storesToCheck_1_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11584.4]
  assign entriesToCheck_1_8 = _T_12856 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11585.4]
  assign _T_12858 = storesToCheck_1_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11586.4]
  assign entriesToCheck_1_9 = _T_12858 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11587.4]
  assign _T_12860 = storesToCheck_1_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11588.4]
  assign entriesToCheck_1_10 = _T_12860 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11589.4]
  assign _T_12862 = storesToCheck_1_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11590.4]
  assign entriesToCheck_1_11 = _T_12862 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11591.4]
  assign _T_12864 = storesToCheck_1_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11592.4]
  assign entriesToCheck_1_12 = _T_12864 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11593.4]
  assign _T_12866 = storesToCheck_1_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11594.4]
  assign entriesToCheck_1_13 = _T_12866 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11595.4]
  assign _T_12868 = storesToCheck_1_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11596.4]
  assign entriesToCheck_1_14 = _T_12868 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11597.4]
  assign _T_12870 = storesToCheck_1_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11598.4]
  assign entriesToCheck_1_15 = _T_12870 & checkBits_1; // @[AxiLoadQueue.scala 140:26:@11599.4]
  assign _T_12872 = storesToCheck_2_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11616.4]
  assign entriesToCheck_2_0 = _T_12872 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11617.4]
  assign _T_12874 = storesToCheck_2_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11618.4]
  assign entriesToCheck_2_1 = _T_12874 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11619.4]
  assign _T_12876 = storesToCheck_2_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11620.4]
  assign entriesToCheck_2_2 = _T_12876 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11621.4]
  assign _T_12878 = storesToCheck_2_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11622.4]
  assign entriesToCheck_2_3 = _T_12878 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11623.4]
  assign _T_12880 = storesToCheck_2_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11624.4]
  assign entriesToCheck_2_4 = _T_12880 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11625.4]
  assign _T_12882 = storesToCheck_2_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11626.4]
  assign entriesToCheck_2_5 = _T_12882 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11627.4]
  assign _T_12884 = storesToCheck_2_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11628.4]
  assign entriesToCheck_2_6 = _T_12884 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11629.4]
  assign _T_12886 = storesToCheck_2_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11630.4]
  assign entriesToCheck_2_7 = _T_12886 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11631.4]
  assign _T_12888 = storesToCheck_2_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11632.4]
  assign entriesToCheck_2_8 = _T_12888 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11633.4]
  assign _T_12890 = storesToCheck_2_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11634.4]
  assign entriesToCheck_2_9 = _T_12890 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11635.4]
  assign _T_12892 = storesToCheck_2_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11636.4]
  assign entriesToCheck_2_10 = _T_12892 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11637.4]
  assign _T_12894 = storesToCheck_2_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11638.4]
  assign entriesToCheck_2_11 = _T_12894 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11639.4]
  assign _T_12896 = storesToCheck_2_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11640.4]
  assign entriesToCheck_2_12 = _T_12896 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11641.4]
  assign _T_12898 = storesToCheck_2_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11642.4]
  assign entriesToCheck_2_13 = _T_12898 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11643.4]
  assign _T_12900 = storesToCheck_2_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11644.4]
  assign entriesToCheck_2_14 = _T_12900 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11645.4]
  assign _T_12902 = storesToCheck_2_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11646.4]
  assign entriesToCheck_2_15 = _T_12902 & checkBits_2; // @[AxiLoadQueue.scala 140:26:@11647.4]
  assign _T_12904 = storesToCheck_3_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11664.4]
  assign entriesToCheck_3_0 = _T_12904 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11665.4]
  assign _T_12906 = storesToCheck_3_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11666.4]
  assign entriesToCheck_3_1 = _T_12906 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11667.4]
  assign _T_12908 = storesToCheck_3_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11668.4]
  assign entriesToCheck_3_2 = _T_12908 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11669.4]
  assign _T_12910 = storesToCheck_3_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11670.4]
  assign entriesToCheck_3_3 = _T_12910 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11671.4]
  assign _T_12912 = storesToCheck_3_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11672.4]
  assign entriesToCheck_3_4 = _T_12912 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11673.4]
  assign _T_12914 = storesToCheck_3_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11674.4]
  assign entriesToCheck_3_5 = _T_12914 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11675.4]
  assign _T_12916 = storesToCheck_3_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11676.4]
  assign entriesToCheck_3_6 = _T_12916 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11677.4]
  assign _T_12918 = storesToCheck_3_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11678.4]
  assign entriesToCheck_3_7 = _T_12918 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11679.4]
  assign _T_12920 = storesToCheck_3_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11680.4]
  assign entriesToCheck_3_8 = _T_12920 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11681.4]
  assign _T_12922 = storesToCheck_3_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11682.4]
  assign entriesToCheck_3_9 = _T_12922 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11683.4]
  assign _T_12924 = storesToCheck_3_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11684.4]
  assign entriesToCheck_3_10 = _T_12924 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11685.4]
  assign _T_12926 = storesToCheck_3_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11686.4]
  assign entriesToCheck_3_11 = _T_12926 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11687.4]
  assign _T_12928 = storesToCheck_3_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11688.4]
  assign entriesToCheck_3_12 = _T_12928 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11689.4]
  assign _T_12930 = storesToCheck_3_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11690.4]
  assign entriesToCheck_3_13 = _T_12930 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11691.4]
  assign _T_12932 = storesToCheck_3_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11692.4]
  assign entriesToCheck_3_14 = _T_12932 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11693.4]
  assign _T_12934 = storesToCheck_3_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11694.4]
  assign entriesToCheck_3_15 = _T_12934 & checkBits_3; // @[AxiLoadQueue.scala 140:26:@11695.4]
  assign _T_12936 = storesToCheck_4_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11712.4]
  assign entriesToCheck_4_0 = _T_12936 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11713.4]
  assign _T_12938 = storesToCheck_4_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11714.4]
  assign entriesToCheck_4_1 = _T_12938 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11715.4]
  assign _T_12940 = storesToCheck_4_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11716.4]
  assign entriesToCheck_4_2 = _T_12940 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11717.4]
  assign _T_12942 = storesToCheck_4_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11718.4]
  assign entriesToCheck_4_3 = _T_12942 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11719.4]
  assign _T_12944 = storesToCheck_4_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11720.4]
  assign entriesToCheck_4_4 = _T_12944 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11721.4]
  assign _T_12946 = storesToCheck_4_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11722.4]
  assign entriesToCheck_4_5 = _T_12946 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11723.4]
  assign _T_12948 = storesToCheck_4_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11724.4]
  assign entriesToCheck_4_6 = _T_12948 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11725.4]
  assign _T_12950 = storesToCheck_4_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11726.4]
  assign entriesToCheck_4_7 = _T_12950 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11727.4]
  assign _T_12952 = storesToCheck_4_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11728.4]
  assign entriesToCheck_4_8 = _T_12952 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11729.4]
  assign _T_12954 = storesToCheck_4_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11730.4]
  assign entriesToCheck_4_9 = _T_12954 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11731.4]
  assign _T_12956 = storesToCheck_4_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11732.4]
  assign entriesToCheck_4_10 = _T_12956 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11733.4]
  assign _T_12958 = storesToCheck_4_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11734.4]
  assign entriesToCheck_4_11 = _T_12958 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11735.4]
  assign _T_12960 = storesToCheck_4_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11736.4]
  assign entriesToCheck_4_12 = _T_12960 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11737.4]
  assign _T_12962 = storesToCheck_4_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11738.4]
  assign entriesToCheck_4_13 = _T_12962 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11739.4]
  assign _T_12964 = storesToCheck_4_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11740.4]
  assign entriesToCheck_4_14 = _T_12964 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11741.4]
  assign _T_12966 = storesToCheck_4_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11742.4]
  assign entriesToCheck_4_15 = _T_12966 & checkBits_4; // @[AxiLoadQueue.scala 140:26:@11743.4]
  assign _T_12968 = storesToCheck_5_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11760.4]
  assign entriesToCheck_5_0 = _T_12968 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11761.4]
  assign _T_12970 = storesToCheck_5_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11762.4]
  assign entriesToCheck_5_1 = _T_12970 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11763.4]
  assign _T_12972 = storesToCheck_5_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11764.4]
  assign entriesToCheck_5_2 = _T_12972 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11765.4]
  assign _T_12974 = storesToCheck_5_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11766.4]
  assign entriesToCheck_5_3 = _T_12974 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11767.4]
  assign _T_12976 = storesToCheck_5_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11768.4]
  assign entriesToCheck_5_4 = _T_12976 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11769.4]
  assign _T_12978 = storesToCheck_5_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11770.4]
  assign entriesToCheck_5_5 = _T_12978 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11771.4]
  assign _T_12980 = storesToCheck_5_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11772.4]
  assign entriesToCheck_5_6 = _T_12980 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11773.4]
  assign _T_12982 = storesToCheck_5_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11774.4]
  assign entriesToCheck_5_7 = _T_12982 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11775.4]
  assign _T_12984 = storesToCheck_5_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11776.4]
  assign entriesToCheck_5_8 = _T_12984 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11777.4]
  assign _T_12986 = storesToCheck_5_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11778.4]
  assign entriesToCheck_5_9 = _T_12986 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11779.4]
  assign _T_12988 = storesToCheck_5_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11780.4]
  assign entriesToCheck_5_10 = _T_12988 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11781.4]
  assign _T_12990 = storesToCheck_5_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11782.4]
  assign entriesToCheck_5_11 = _T_12990 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11783.4]
  assign _T_12992 = storesToCheck_5_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11784.4]
  assign entriesToCheck_5_12 = _T_12992 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11785.4]
  assign _T_12994 = storesToCheck_5_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11786.4]
  assign entriesToCheck_5_13 = _T_12994 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11787.4]
  assign _T_12996 = storesToCheck_5_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11788.4]
  assign entriesToCheck_5_14 = _T_12996 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11789.4]
  assign _T_12998 = storesToCheck_5_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11790.4]
  assign entriesToCheck_5_15 = _T_12998 & checkBits_5; // @[AxiLoadQueue.scala 140:26:@11791.4]
  assign _T_13000 = storesToCheck_6_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11808.4]
  assign entriesToCheck_6_0 = _T_13000 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11809.4]
  assign _T_13002 = storesToCheck_6_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11810.4]
  assign entriesToCheck_6_1 = _T_13002 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11811.4]
  assign _T_13004 = storesToCheck_6_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11812.4]
  assign entriesToCheck_6_2 = _T_13004 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11813.4]
  assign _T_13006 = storesToCheck_6_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11814.4]
  assign entriesToCheck_6_3 = _T_13006 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11815.4]
  assign _T_13008 = storesToCheck_6_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11816.4]
  assign entriesToCheck_6_4 = _T_13008 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11817.4]
  assign _T_13010 = storesToCheck_6_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11818.4]
  assign entriesToCheck_6_5 = _T_13010 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11819.4]
  assign _T_13012 = storesToCheck_6_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11820.4]
  assign entriesToCheck_6_6 = _T_13012 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11821.4]
  assign _T_13014 = storesToCheck_6_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11822.4]
  assign entriesToCheck_6_7 = _T_13014 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11823.4]
  assign _T_13016 = storesToCheck_6_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11824.4]
  assign entriesToCheck_6_8 = _T_13016 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11825.4]
  assign _T_13018 = storesToCheck_6_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11826.4]
  assign entriesToCheck_6_9 = _T_13018 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11827.4]
  assign _T_13020 = storesToCheck_6_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11828.4]
  assign entriesToCheck_6_10 = _T_13020 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11829.4]
  assign _T_13022 = storesToCheck_6_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11830.4]
  assign entriesToCheck_6_11 = _T_13022 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11831.4]
  assign _T_13024 = storesToCheck_6_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11832.4]
  assign entriesToCheck_6_12 = _T_13024 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11833.4]
  assign _T_13026 = storesToCheck_6_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11834.4]
  assign entriesToCheck_6_13 = _T_13026 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11835.4]
  assign _T_13028 = storesToCheck_6_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11836.4]
  assign entriesToCheck_6_14 = _T_13028 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11837.4]
  assign _T_13030 = storesToCheck_6_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11838.4]
  assign entriesToCheck_6_15 = _T_13030 & checkBits_6; // @[AxiLoadQueue.scala 140:26:@11839.4]
  assign _T_13032 = storesToCheck_7_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11856.4]
  assign entriesToCheck_7_0 = _T_13032 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11857.4]
  assign _T_13034 = storesToCheck_7_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11858.4]
  assign entriesToCheck_7_1 = _T_13034 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11859.4]
  assign _T_13036 = storesToCheck_7_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11860.4]
  assign entriesToCheck_7_2 = _T_13036 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11861.4]
  assign _T_13038 = storesToCheck_7_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11862.4]
  assign entriesToCheck_7_3 = _T_13038 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11863.4]
  assign _T_13040 = storesToCheck_7_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11864.4]
  assign entriesToCheck_7_4 = _T_13040 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11865.4]
  assign _T_13042 = storesToCheck_7_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11866.4]
  assign entriesToCheck_7_5 = _T_13042 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11867.4]
  assign _T_13044 = storesToCheck_7_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11868.4]
  assign entriesToCheck_7_6 = _T_13044 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11869.4]
  assign _T_13046 = storesToCheck_7_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11870.4]
  assign entriesToCheck_7_7 = _T_13046 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11871.4]
  assign _T_13048 = storesToCheck_7_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11872.4]
  assign entriesToCheck_7_8 = _T_13048 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11873.4]
  assign _T_13050 = storesToCheck_7_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11874.4]
  assign entriesToCheck_7_9 = _T_13050 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11875.4]
  assign _T_13052 = storesToCheck_7_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11876.4]
  assign entriesToCheck_7_10 = _T_13052 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11877.4]
  assign _T_13054 = storesToCheck_7_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11878.4]
  assign entriesToCheck_7_11 = _T_13054 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11879.4]
  assign _T_13056 = storesToCheck_7_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11880.4]
  assign entriesToCheck_7_12 = _T_13056 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11881.4]
  assign _T_13058 = storesToCheck_7_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11882.4]
  assign entriesToCheck_7_13 = _T_13058 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11883.4]
  assign _T_13060 = storesToCheck_7_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11884.4]
  assign entriesToCheck_7_14 = _T_13060 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11885.4]
  assign _T_13062 = storesToCheck_7_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11886.4]
  assign entriesToCheck_7_15 = _T_13062 & checkBits_7; // @[AxiLoadQueue.scala 140:26:@11887.4]
  assign _T_13064 = storesToCheck_8_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11904.4]
  assign entriesToCheck_8_0 = _T_13064 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11905.4]
  assign _T_13066 = storesToCheck_8_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11906.4]
  assign entriesToCheck_8_1 = _T_13066 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11907.4]
  assign _T_13068 = storesToCheck_8_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11908.4]
  assign entriesToCheck_8_2 = _T_13068 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11909.4]
  assign _T_13070 = storesToCheck_8_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11910.4]
  assign entriesToCheck_8_3 = _T_13070 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11911.4]
  assign _T_13072 = storesToCheck_8_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11912.4]
  assign entriesToCheck_8_4 = _T_13072 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11913.4]
  assign _T_13074 = storesToCheck_8_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11914.4]
  assign entriesToCheck_8_5 = _T_13074 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11915.4]
  assign _T_13076 = storesToCheck_8_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11916.4]
  assign entriesToCheck_8_6 = _T_13076 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11917.4]
  assign _T_13078 = storesToCheck_8_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11918.4]
  assign entriesToCheck_8_7 = _T_13078 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11919.4]
  assign _T_13080 = storesToCheck_8_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11920.4]
  assign entriesToCheck_8_8 = _T_13080 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11921.4]
  assign _T_13082 = storesToCheck_8_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11922.4]
  assign entriesToCheck_8_9 = _T_13082 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11923.4]
  assign _T_13084 = storesToCheck_8_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11924.4]
  assign entriesToCheck_8_10 = _T_13084 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11925.4]
  assign _T_13086 = storesToCheck_8_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11926.4]
  assign entriesToCheck_8_11 = _T_13086 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11927.4]
  assign _T_13088 = storesToCheck_8_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11928.4]
  assign entriesToCheck_8_12 = _T_13088 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11929.4]
  assign _T_13090 = storesToCheck_8_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11930.4]
  assign entriesToCheck_8_13 = _T_13090 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11931.4]
  assign _T_13092 = storesToCheck_8_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11932.4]
  assign entriesToCheck_8_14 = _T_13092 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11933.4]
  assign _T_13094 = storesToCheck_8_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11934.4]
  assign entriesToCheck_8_15 = _T_13094 & checkBits_8; // @[AxiLoadQueue.scala 140:26:@11935.4]
  assign _T_13096 = storesToCheck_9_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@11952.4]
  assign entriesToCheck_9_0 = _T_13096 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11953.4]
  assign _T_13098 = storesToCheck_9_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@11954.4]
  assign entriesToCheck_9_1 = _T_13098 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11955.4]
  assign _T_13100 = storesToCheck_9_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@11956.4]
  assign entriesToCheck_9_2 = _T_13100 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11957.4]
  assign _T_13102 = storesToCheck_9_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@11958.4]
  assign entriesToCheck_9_3 = _T_13102 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11959.4]
  assign _T_13104 = storesToCheck_9_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@11960.4]
  assign entriesToCheck_9_4 = _T_13104 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11961.4]
  assign _T_13106 = storesToCheck_9_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@11962.4]
  assign entriesToCheck_9_5 = _T_13106 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11963.4]
  assign _T_13108 = storesToCheck_9_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@11964.4]
  assign entriesToCheck_9_6 = _T_13108 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11965.4]
  assign _T_13110 = storesToCheck_9_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@11966.4]
  assign entriesToCheck_9_7 = _T_13110 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11967.4]
  assign _T_13112 = storesToCheck_9_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@11968.4]
  assign entriesToCheck_9_8 = _T_13112 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11969.4]
  assign _T_13114 = storesToCheck_9_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@11970.4]
  assign entriesToCheck_9_9 = _T_13114 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11971.4]
  assign _T_13116 = storesToCheck_9_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@11972.4]
  assign entriesToCheck_9_10 = _T_13116 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11973.4]
  assign _T_13118 = storesToCheck_9_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@11974.4]
  assign entriesToCheck_9_11 = _T_13118 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11975.4]
  assign _T_13120 = storesToCheck_9_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@11976.4]
  assign entriesToCheck_9_12 = _T_13120 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11977.4]
  assign _T_13122 = storesToCheck_9_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@11978.4]
  assign entriesToCheck_9_13 = _T_13122 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11979.4]
  assign _T_13124 = storesToCheck_9_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@11980.4]
  assign entriesToCheck_9_14 = _T_13124 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11981.4]
  assign _T_13126 = storesToCheck_9_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@11982.4]
  assign entriesToCheck_9_15 = _T_13126 & checkBits_9; // @[AxiLoadQueue.scala 140:26:@11983.4]
  assign _T_13128 = storesToCheck_10_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@12000.4]
  assign entriesToCheck_10_0 = _T_13128 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12001.4]
  assign _T_13130 = storesToCheck_10_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@12002.4]
  assign entriesToCheck_10_1 = _T_13130 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12003.4]
  assign _T_13132 = storesToCheck_10_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@12004.4]
  assign entriesToCheck_10_2 = _T_13132 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12005.4]
  assign _T_13134 = storesToCheck_10_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@12006.4]
  assign entriesToCheck_10_3 = _T_13134 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12007.4]
  assign _T_13136 = storesToCheck_10_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@12008.4]
  assign entriesToCheck_10_4 = _T_13136 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12009.4]
  assign _T_13138 = storesToCheck_10_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@12010.4]
  assign entriesToCheck_10_5 = _T_13138 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12011.4]
  assign _T_13140 = storesToCheck_10_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@12012.4]
  assign entriesToCheck_10_6 = _T_13140 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12013.4]
  assign _T_13142 = storesToCheck_10_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@12014.4]
  assign entriesToCheck_10_7 = _T_13142 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12015.4]
  assign _T_13144 = storesToCheck_10_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@12016.4]
  assign entriesToCheck_10_8 = _T_13144 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12017.4]
  assign _T_13146 = storesToCheck_10_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@12018.4]
  assign entriesToCheck_10_9 = _T_13146 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12019.4]
  assign _T_13148 = storesToCheck_10_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@12020.4]
  assign entriesToCheck_10_10 = _T_13148 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12021.4]
  assign _T_13150 = storesToCheck_10_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@12022.4]
  assign entriesToCheck_10_11 = _T_13150 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12023.4]
  assign _T_13152 = storesToCheck_10_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@12024.4]
  assign entriesToCheck_10_12 = _T_13152 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12025.4]
  assign _T_13154 = storesToCheck_10_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@12026.4]
  assign entriesToCheck_10_13 = _T_13154 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12027.4]
  assign _T_13156 = storesToCheck_10_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@12028.4]
  assign entriesToCheck_10_14 = _T_13156 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12029.4]
  assign _T_13158 = storesToCheck_10_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@12030.4]
  assign entriesToCheck_10_15 = _T_13158 & checkBits_10; // @[AxiLoadQueue.scala 140:26:@12031.4]
  assign _T_13160 = storesToCheck_11_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@12048.4]
  assign entriesToCheck_11_0 = _T_13160 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12049.4]
  assign _T_13162 = storesToCheck_11_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@12050.4]
  assign entriesToCheck_11_1 = _T_13162 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12051.4]
  assign _T_13164 = storesToCheck_11_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@12052.4]
  assign entriesToCheck_11_2 = _T_13164 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12053.4]
  assign _T_13166 = storesToCheck_11_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@12054.4]
  assign entriesToCheck_11_3 = _T_13166 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12055.4]
  assign _T_13168 = storesToCheck_11_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@12056.4]
  assign entriesToCheck_11_4 = _T_13168 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12057.4]
  assign _T_13170 = storesToCheck_11_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@12058.4]
  assign entriesToCheck_11_5 = _T_13170 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12059.4]
  assign _T_13172 = storesToCheck_11_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@12060.4]
  assign entriesToCheck_11_6 = _T_13172 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12061.4]
  assign _T_13174 = storesToCheck_11_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@12062.4]
  assign entriesToCheck_11_7 = _T_13174 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12063.4]
  assign _T_13176 = storesToCheck_11_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@12064.4]
  assign entriesToCheck_11_8 = _T_13176 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12065.4]
  assign _T_13178 = storesToCheck_11_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@12066.4]
  assign entriesToCheck_11_9 = _T_13178 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12067.4]
  assign _T_13180 = storesToCheck_11_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@12068.4]
  assign entriesToCheck_11_10 = _T_13180 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12069.4]
  assign _T_13182 = storesToCheck_11_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@12070.4]
  assign entriesToCheck_11_11 = _T_13182 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12071.4]
  assign _T_13184 = storesToCheck_11_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@12072.4]
  assign entriesToCheck_11_12 = _T_13184 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12073.4]
  assign _T_13186 = storesToCheck_11_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@12074.4]
  assign entriesToCheck_11_13 = _T_13186 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12075.4]
  assign _T_13188 = storesToCheck_11_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@12076.4]
  assign entriesToCheck_11_14 = _T_13188 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12077.4]
  assign _T_13190 = storesToCheck_11_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@12078.4]
  assign entriesToCheck_11_15 = _T_13190 & checkBits_11; // @[AxiLoadQueue.scala 140:26:@12079.4]
  assign _T_13192 = storesToCheck_12_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@12096.4]
  assign entriesToCheck_12_0 = _T_13192 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12097.4]
  assign _T_13194 = storesToCheck_12_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@12098.4]
  assign entriesToCheck_12_1 = _T_13194 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12099.4]
  assign _T_13196 = storesToCheck_12_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@12100.4]
  assign entriesToCheck_12_2 = _T_13196 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12101.4]
  assign _T_13198 = storesToCheck_12_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@12102.4]
  assign entriesToCheck_12_3 = _T_13198 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12103.4]
  assign _T_13200 = storesToCheck_12_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@12104.4]
  assign entriesToCheck_12_4 = _T_13200 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12105.4]
  assign _T_13202 = storesToCheck_12_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@12106.4]
  assign entriesToCheck_12_5 = _T_13202 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12107.4]
  assign _T_13204 = storesToCheck_12_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@12108.4]
  assign entriesToCheck_12_6 = _T_13204 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12109.4]
  assign _T_13206 = storesToCheck_12_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@12110.4]
  assign entriesToCheck_12_7 = _T_13206 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12111.4]
  assign _T_13208 = storesToCheck_12_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@12112.4]
  assign entriesToCheck_12_8 = _T_13208 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12113.4]
  assign _T_13210 = storesToCheck_12_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@12114.4]
  assign entriesToCheck_12_9 = _T_13210 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12115.4]
  assign _T_13212 = storesToCheck_12_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@12116.4]
  assign entriesToCheck_12_10 = _T_13212 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12117.4]
  assign _T_13214 = storesToCheck_12_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@12118.4]
  assign entriesToCheck_12_11 = _T_13214 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12119.4]
  assign _T_13216 = storesToCheck_12_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@12120.4]
  assign entriesToCheck_12_12 = _T_13216 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12121.4]
  assign _T_13218 = storesToCheck_12_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@12122.4]
  assign entriesToCheck_12_13 = _T_13218 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12123.4]
  assign _T_13220 = storesToCheck_12_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@12124.4]
  assign entriesToCheck_12_14 = _T_13220 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12125.4]
  assign _T_13222 = storesToCheck_12_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@12126.4]
  assign entriesToCheck_12_15 = _T_13222 & checkBits_12; // @[AxiLoadQueue.scala 140:26:@12127.4]
  assign _T_13224 = storesToCheck_13_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@12144.4]
  assign entriesToCheck_13_0 = _T_13224 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12145.4]
  assign _T_13226 = storesToCheck_13_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@12146.4]
  assign entriesToCheck_13_1 = _T_13226 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12147.4]
  assign _T_13228 = storesToCheck_13_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@12148.4]
  assign entriesToCheck_13_2 = _T_13228 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12149.4]
  assign _T_13230 = storesToCheck_13_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@12150.4]
  assign entriesToCheck_13_3 = _T_13230 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12151.4]
  assign _T_13232 = storesToCheck_13_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@12152.4]
  assign entriesToCheck_13_4 = _T_13232 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12153.4]
  assign _T_13234 = storesToCheck_13_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@12154.4]
  assign entriesToCheck_13_5 = _T_13234 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12155.4]
  assign _T_13236 = storesToCheck_13_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@12156.4]
  assign entriesToCheck_13_6 = _T_13236 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12157.4]
  assign _T_13238 = storesToCheck_13_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@12158.4]
  assign entriesToCheck_13_7 = _T_13238 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12159.4]
  assign _T_13240 = storesToCheck_13_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@12160.4]
  assign entriesToCheck_13_8 = _T_13240 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12161.4]
  assign _T_13242 = storesToCheck_13_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@12162.4]
  assign entriesToCheck_13_9 = _T_13242 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12163.4]
  assign _T_13244 = storesToCheck_13_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@12164.4]
  assign entriesToCheck_13_10 = _T_13244 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12165.4]
  assign _T_13246 = storesToCheck_13_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@12166.4]
  assign entriesToCheck_13_11 = _T_13246 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12167.4]
  assign _T_13248 = storesToCheck_13_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@12168.4]
  assign entriesToCheck_13_12 = _T_13248 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12169.4]
  assign _T_13250 = storesToCheck_13_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@12170.4]
  assign entriesToCheck_13_13 = _T_13250 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12171.4]
  assign _T_13252 = storesToCheck_13_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@12172.4]
  assign entriesToCheck_13_14 = _T_13252 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12173.4]
  assign _T_13254 = storesToCheck_13_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@12174.4]
  assign entriesToCheck_13_15 = _T_13254 & checkBits_13; // @[AxiLoadQueue.scala 140:26:@12175.4]
  assign _T_13256 = storesToCheck_14_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@12192.4]
  assign entriesToCheck_14_0 = _T_13256 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12193.4]
  assign _T_13258 = storesToCheck_14_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@12194.4]
  assign entriesToCheck_14_1 = _T_13258 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12195.4]
  assign _T_13260 = storesToCheck_14_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@12196.4]
  assign entriesToCheck_14_2 = _T_13260 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12197.4]
  assign _T_13262 = storesToCheck_14_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@12198.4]
  assign entriesToCheck_14_3 = _T_13262 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12199.4]
  assign _T_13264 = storesToCheck_14_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@12200.4]
  assign entriesToCheck_14_4 = _T_13264 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12201.4]
  assign _T_13266 = storesToCheck_14_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@12202.4]
  assign entriesToCheck_14_5 = _T_13266 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12203.4]
  assign _T_13268 = storesToCheck_14_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@12204.4]
  assign entriesToCheck_14_6 = _T_13268 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12205.4]
  assign _T_13270 = storesToCheck_14_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@12206.4]
  assign entriesToCheck_14_7 = _T_13270 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12207.4]
  assign _T_13272 = storesToCheck_14_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@12208.4]
  assign entriesToCheck_14_8 = _T_13272 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12209.4]
  assign _T_13274 = storesToCheck_14_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@12210.4]
  assign entriesToCheck_14_9 = _T_13274 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12211.4]
  assign _T_13276 = storesToCheck_14_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@12212.4]
  assign entriesToCheck_14_10 = _T_13276 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12213.4]
  assign _T_13278 = storesToCheck_14_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@12214.4]
  assign entriesToCheck_14_11 = _T_13278 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12215.4]
  assign _T_13280 = storesToCheck_14_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@12216.4]
  assign entriesToCheck_14_12 = _T_13280 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12217.4]
  assign _T_13282 = storesToCheck_14_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@12218.4]
  assign entriesToCheck_14_13 = _T_13282 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12219.4]
  assign _T_13284 = storesToCheck_14_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@12220.4]
  assign entriesToCheck_14_14 = _T_13284 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12221.4]
  assign _T_13286 = storesToCheck_14_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@12222.4]
  assign entriesToCheck_14_15 = _T_13286 & checkBits_14; // @[AxiLoadQueue.scala 140:26:@12223.4]
  assign _T_13288 = storesToCheck_15_0 & validEntriesInStoreQ_0; // @[AxiLoadQueue.scala 140:18:@12240.4]
  assign entriesToCheck_15_0 = _T_13288 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12241.4]
  assign _T_13290 = storesToCheck_15_1 & validEntriesInStoreQ_1; // @[AxiLoadQueue.scala 140:18:@12242.4]
  assign entriesToCheck_15_1 = _T_13290 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12243.4]
  assign _T_13292 = storesToCheck_15_2 & validEntriesInStoreQ_2; // @[AxiLoadQueue.scala 140:18:@12244.4]
  assign entriesToCheck_15_2 = _T_13292 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12245.4]
  assign _T_13294 = storesToCheck_15_3 & validEntriesInStoreQ_3; // @[AxiLoadQueue.scala 140:18:@12246.4]
  assign entriesToCheck_15_3 = _T_13294 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12247.4]
  assign _T_13296 = storesToCheck_15_4 & validEntriesInStoreQ_4; // @[AxiLoadQueue.scala 140:18:@12248.4]
  assign entriesToCheck_15_4 = _T_13296 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12249.4]
  assign _T_13298 = storesToCheck_15_5 & validEntriesInStoreQ_5; // @[AxiLoadQueue.scala 140:18:@12250.4]
  assign entriesToCheck_15_5 = _T_13298 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12251.4]
  assign _T_13300 = storesToCheck_15_6 & validEntriesInStoreQ_6; // @[AxiLoadQueue.scala 140:18:@12252.4]
  assign entriesToCheck_15_6 = _T_13300 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12253.4]
  assign _T_13302 = storesToCheck_15_7 & validEntriesInStoreQ_7; // @[AxiLoadQueue.scala 140:18:@12254.4]
  assign entriesToCheck_15_7 = _T_13302 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12255.4]
  assign _T_13304 = storesToCheck_15_8 & validEntriesInStoreQ_8; // @[AxiLoadQueue.scala 140:18:@12256.4]
  assign entriesToCheck_15_8 = _T_13304 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12257.4]
  assign _T_13306 = storesToCheck_15_9 & validEntriesInStoreQ_9; // @[AxiLoadQueue.scala 140:18:@12258.4]
  assign entriesToCheck_15_9 = _T_13306 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12259.4]
  assign _T_13308 = storesToCheck_15_10 & validEntriesInStoreQ_10; // @[AxiLoadQueue.scala 140:18:@12260.4]
  assign entriesToCheck_15_10 = _T_13308 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12261.4]
  assign _T_13310 = storesToCheck_15_11 & validEntriesInStoreQ_11; // @[AxiLoadQueue.scala 140:18:@12262.4]
  assign entriesToCheck_15_11 = _T_13310 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12263.4]
  assign _T_13312 = storesToCheck_15_12 & validEntriesInStoreQ_12; // @[AxiLoadQueue.scala 140:18:@12264.4]
  assign entriesToCheck_15_12 = _T_13312 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12265.4]
  assign _T_13314 = storesToCheck_15_13 & validEntriesInStoreQ_13; // @[AxiLoadQueue.scala 140:18:@12266.4]
  assign entriesToCheck_15_13 = _T_13314 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12267.4]
  assign _T_13316 = storesToCheck_15_14 & validEntriesInStoreQ_14; // @[AxiLoadQueue.scala 140:18:@12268.4]
  assign entriesToCheck_15_14 = _T_13316 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12269.4]
  assign _T_13318 = storesToCheck_15_15 & validEntriesInStoreQ_15; // @[AxiLoadQueue.scala 140:18:@12270.4]
  assign entriesToCheck_15_15 = _T_13318 & checkBits_15; // @[AxiLoadQueue.scala 140:26:@12271.4]
  assign _T_14550 = entriesToCheck_0_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12289.4]
  assign _T_14551 = _T_14550 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12290.4]
  assign _T_14552 = addrQ_0 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12291.4]
  assign conflict_0_0 = _T_14551 & _T_14552; // @[AxiLoadQueue.scala 151:68:@12292.4]
  assign _T_14554 = entriesToCheck_0_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12294.4]
  assign _T_14555 = _T_14554 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12295.4]
  assign _T_14556 = addrQ_0 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12296.4]
  assign conflict_0_1 = _T_14555 & _T_14556; // @[AxiLoadQueue.scala 151:68:@12297.4]
  assign _T_14558 = entriesToCheck_0_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12299.4]
  assign _T_14559 = _T_14558 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12300.4]
  assign _T_14560 = addrQ_0 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12301.4]
  assign conflict_0_2 = _T_14559 & _T_14560; // @[AxiLoadQueue.scala 151:68:@12302.4]
  assign _T_14562 = entriesToCheck_0_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12304.4]
  assign _T_14563 = _T_14562 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12305.4]
  assign _T_14564 = addrQ_0 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12306.4]
  assign conflict_0_3 = _T_14563 & _T_14564; // @[AxiLoadQueue.scala 151:68:@12307.4]
  assign _T_14566 = entriesToCheck_0_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12309.4]
  assign _T_14567 = _T_14566 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12310.4]
  assign _T_14568 = addrQ_0 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12311.4]
  assign conflict_0_4 = _T_14567 & _T_14568; // @[AxiLoadQueue.scala 151:68:@12312.4]
  assign _T_14570 = entriesToCheck_0_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12314.4]
  assign _T_14571 = _T_14570 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12315.4]
  assign _T_14572 = addrQ_0 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12316.4]
  assign conflict_0_5 = _T_14571 & _T_14572; // @[AxiLoadQueue.scala 151:68:@12317.4]
  assign _T_14574 = entriesToCheck_0_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12319.4]
  assign _T_14575 = _T_14574 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12320.4]
  assign _T_14576 = addrQ_0 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12321.4]
  assign conflict_0_6 = _T_14575 & _T_14576; // @[AxiLoadQueue.scala 151:68:@12322.4]
  assign _T_14578 = entriesToCheck_0_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12324.4]
  assign _T_14579 = _T_14578 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12325.4]
  assign _T_14580 = addrQ_0 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12326.4]
  assign conflict_0_7 = _T_14579 & _T_14580; // @[AxiLoadQueue.scala 151:68:@12327.4]
  assign _T_14582 = entriesToCheck_0_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12329.4]
  assign _T_14583 = _T_14582 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12330.4]
  assign _T_14584 = addrQ_0 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12331.4]
  assign conflict_0_8 = _T_14583 & _T_14584; // @[AxiLoadQueue.scala 151:68:@12332.4]
  assign _T_14586 = entriesToCheck_0_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12334.4]
  assign _T_14587 = _T_14586 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12335.4]
  assign _T_14588 = addrQ_0 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12336.4]
  assign conflict_0_9 = _T_14587 & _T_14588; // @[AxiLoadQueue.scala 151:68:@12337.4]
  assign _T_14590 = entriesToCheck_0_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12339.4]
  assign _T_14591 = _T_14590 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12340.4]
  assign _T_14592 = addrQ_0 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12341.4]
  assign conflict_0_10 = _T_14591 & _T_14592; // @[AxiLoadQueue.scala 151:68:@12342.4]
  assign _T_14594 = entriesToCheck_0_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12344.4]
  assign _T_14595 = _T_14594 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12345.4]
  assign _T_14596 = addrQ_0 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12346.4]
  assign conflict_0_11 = _T_14595 & _T_14596; // @[AxiLoadQueue.scala 151:68:@12347.4]
  assign _T_14598 = entriesToCheck_0_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12349.4]
  assign _T_14599 = _T_14598 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12350.4]
  assign _T_14600 = addrQ_0 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12351.4]
  assign conflict_0_12 = _T_14599 & _T_14600; // @[AxiLoadQueue.scala 151:68:@12352.4]
  assign _T_14602 = entriesToCheck_0_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12354.4]
  assign _T_14603 = _T_14602 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12355.4]
  assign _T_14604 = addrQ_0 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12356.4]
  assign conflict_0_13 = _T_14603 & _T_14604; // @[AxiLoadQueue.scala 151:68:@12357.4]
  assign _T_14606 = entriesToCheck_0_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12359.4]
  assign _T_14607 = _T_14606 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12360.4]
  assign _T_14608 = addrQ_0 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12361.4]
  assign conflict_0_14 = _T_14607 & _T_14608; // @[AxiLoadQueue.scala 151:68:@12362.4]
  assign _T_14610 = entriesToCheck_0_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12364.4]
  assign _T_14611 = _T_14610 & addrKnown_0; // @[AxiLoadQueue.scala 151:41:@12365.4]
  assign _T_14612 = addrQ_0 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12366.4]
  assign conflict_0_15 = _T_14611 & _T_14612; // @[AxiLoadQueue.scala 151:68:@12367.4]
  assign _T_14614 = entriesToCheck_1_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12369.4]
  assign _T_14615 = _T_14614 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12370.4]
  assign _T_14616 = addrQ_1 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12371.4]
  assign conflict_1_0 = _T_14615 & _T_14616; // @[AxiLoadQueue.scala 151:68:@12372.4]
  assign _T_14618 = entriesToCheck_1_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12374.4]
  assign _T_14619 = _T_14618 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12375.4]
  assign _T_14620 = addrQ_1 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12376.4]
  assign conflict_1_1 = _T_14619 & _T_14620; // @[AxiLoadQueue.scala 151:68:@12377.4]
  assign _T_14622 = entriesToCheck_1_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12379.4]
  assign _T_14623 = _T_14622 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12380.4]
  assign _T_14624 = addrQ_1 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12381.4]
  assign conflict_1_2 = _T_14623 & _T_14624; // @[AxiLoadQueue.scala 151:68:@12382.4]
  assign _T_14626 = entriesToCheck_1_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12384.4]
  assign _T_14627 = _T_14626 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12385.4]
  assign _T_14628 = addrQ_1 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12386.4]
  assign conflict_1_3 = _T_14627 & _T_14628; // @[AxiLoadQueue.scala 151:68:@12387.4]
  assign _T_14630 = entriesToCheck_1_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12389.4]
  assign _T_14631 = _T_14630 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12390.4]
  assign _T_14632 = addrQ_1 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12391.4]
  assign conflict_1_4 = _T_14631 & _T_14632; // @[AxiLoadQueue.scala 151:68:@12392.4]
  assign _T_14634 = entriesToCheck_1_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12394.4]
  assign _T_14635 = _T_14634 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12395.4]
  assign _T_14636 = addrQ_1 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12396.4]
  assign conflict_1_5 = _T_14635 & _T_14636; // @[AxiLoadQueue.scala 151:68:@12397.4]
  assign _T_14638 = entriesToCheck_1_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12399.4]
  assign _T_14639 = _T_14638 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12400.4]
  assign _T_14640 = addrQ_1 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12401.4]
  assign conflict_1_6 = _T_14639 & _T_14640; // @[AxiLoadQueue.scala 151:68:@12402.4]
  assign _T_14642 = entriesToCheck_1_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12404.4]
  assign _T_14643 = _T_14642 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12405.4]
  assign _T_14644 = addrQ_1 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12406.4]
  assign conflict_1_7 = _T_14643 & _T_14644; // @[AxiLoadQueue.scala 151:68:@12407.4]
  assign _T_14646 = entriesToCheck_1_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12409.4]
  assign _T_14647 = _T_14646 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12410.4]
  assign _T_14648 = addrQ_1 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12411.4]
  assign conflict_1_8 = _T_14647 & _T_14648; // @[AxiLoadQueue.scala 151:68:@12412.4]
  assign _T_14650 = entriesToCheck_1_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12414.4]
  assign _T_14651 = _T_14650 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12415.4]
  assign _T_14652 = addrQ_1 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12416.4]
  assign conflict_1_9 = _T_14651 & _T_14652; // @[AxiLoadQueue.scala 151:68:@12417.4]
  assign _T_14654 = entriesToCheck_1_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12419.4]
  assign _T_14655 = _T_14654 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12420.4]
  assign _T_14656 = addrQ_1 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12421.4]
  assign conflict_1_10 = _T_14655 & _T_14656; // @[AxiLoadQueue.scala 151:68:@12422.4]
  assign _T_14658 = entriesToCheck_1_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12424.4]
  assign _T_14659 = _T_14658 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12425.4]
  assign _T_14660 = addrQ_1 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12426.4]
  assign conflict_1_11 = _T_14659 & _T_14660; // @[AxiLoadQueue.scala 151:68:@12427.4]
  assign _T_14662 = entriesToCheck_1_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12429.4]
  assign _T_14663 = _T_14662 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12430.4]
  assign _T_14664 = addrQ_1 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12431.4]
  assign conflict_1_12 = _T_14663 & _T_14664; // @[AxiLoadQueue.scala 151:68:@12432.4]
  assign _T_14666 = entriesToCheck_1_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12434.4]
  assign _T_14667 = _T_14666 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12435.4]
  assign _T_14668 = addrQ_1 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12436.4]
  assign conflict_1_13 = _T_14667 & _T_14668; // @[AxiLoadQueue.scala 151:68:@12437.4]
  assign _T_14670 = entriesToCheck_1_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12439.4]
  assign _T_14671 = _T_14670 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12440.4]
  assign _T_14672 = addrQ_1 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12441.4]
  assign conflict_1_14 = _T_14671 & _T_14672; // @[AxiLoadQueue.scala 151:68:@12442.4]
  assign _T_14674 = entriesToCheck_1_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12444.4]
  assign _T_14675 = _T_14674 & addrKnown_1; // @[AxiLoadQueue.scala 151:41:@12445.4]
  assign _T_14676 = addrQ_1 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12446.4]
  assign conflict_1_15 = _T_14675 & _T_14676; // @[AxiLoadQueue.scala 151:68:@12447.4]
  assign _T_14678 = entriesToCheck_2_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12449.4]
  assign _T_14679 = _T_14678 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12450.4]
  assign _T_14680 = addrQ_2 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12451.4]
  assign conflict_2_0 = _T_14679 & _T_14680; // @[AxiLoadQueue.scala 151:68:@12452.4]
  assign _T_14682 = entriesToCheck_2_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12454.4]
  assign _T_14683 = _T_14682 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12455.4]
  assign _T_14684 = addrQ_2 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12456.4]
  assign conflict_2_1 = _T_14683 & _T_14684; // @[AxiLoadQueue.scala 151:68:@12457.4]
  assign _T_14686 = entriesToCheck_2_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12459.4]
  assign _T_14687 = _T_14686 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12460.4]
  assign _T_14688 = addrQ_2 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12461.4]
  assign conflict_2_2 = _T_14687 & _T_14688; // @[AxiLoadQueue.scala 151:68:@12462.4]
  assign _T_14690 = entriesToCheck_2_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12464.4]
  assign _T_14691 = _T_14690 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12465.4]
  assign _T_14692 = addrQ_2 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12466.4]
  assign conflict_2_3 = _T_14691 & _T_14692; // @[AxiLoadQueue.scala 151:68:@12467.4]
  assign _T_14694 = entriesToCheck_2_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12469.4]
  assign _T_14695 = _T_14694 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12470.4]
  assign _T_14696 = addrQ_2 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12471.4]
  assign conflict_2_4 = _T_14695 & _T_14696; // @[AxiLoadQueue.scala 151:68:@12472.4]
  assign _T_14698 = entriesToCheck_2_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12474.4]
  assign _T_14699 = _T_14698 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12475.4]
  assign _T_14700 = addrQ_2 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12476.4]
  assign conflict_2_5 = _T_14699 & _T_14700; // @[AxiLoadQueue.scala 151:68:@12477.4]
  assign _T_14702 = entriesToCheck_2_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12479.4]
  assign _T_14703 = _T_14702 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12480.4]
  assign _T_14704 = addrQ_2 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12481.4]
  assign conflict_2_6 = _T_14703 & _T_14704; // @[AxiLoadQueue.scala 151:68:@12482.4]
  assign _T_14706 = entriesToCheck_2_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12484.4]
  assign _T_14707 = _T_14706 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12485.4]
  assign _T_14708 = addrQ_2 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12486.4]
  assign conflict_2_7 = _T_14707 & _T_14708; // @[AxiLoadQueue.scala 151:68:@12487.4]
  assign _T_14710 = entriesToCheck_2_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12489.4]
  assign _T_14711 = _T_14710 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12490.4]
  assign _T_14712 = addrQ_2 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12491.4]
  assign conflict_2_8 = _T_14711 & _T_14712; // @[AxiLoadQueue.scala 151:68:@12492.4]
  assign _T_14714 = entriesToCheck_2_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12494.4]
  assign _T_14715 = _T_14714 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12495.4]
  assign _T_14716 = addrQ_2 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12496.4]
  assign conflict_2_9 = _T_14715 & _T_14716; // @[AxiLoadQueue.scala 151:68:@12497.4]
  assign _T_14718 = entriesToCheck_2_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12499.4]
  assign _T_14719 = _T_14718 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12500.4]
  assign _T_14720 = addrQ_2 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12501.4]
  assign conflict_2_10 = _T_14719 & _T_14720; // @[AxiLoadQueue.scala 151:68:@12502.4]
  assign _T_14722 = entriesToCheck_2_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12504.4]
  assign _T_14723 = _T_14722 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12505.4]
  assign _T_14724 = addrQ_2 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12506.4]
  assign conflict_2_11 = _T_14723 & _T_14724; // @[AxiLoadQueue.scala 151:68:@12507.4]
  assign _T_14726 = entriesToCheck_2_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12509.4]
  assign _T_14727 = _T_14726 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12510.4]
  assign _T_14728 = addrQ_2 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12511.4]
  assign conflict_2_12 = _T_14727 & _T_14728; // @[AxiLoadQueue.scala 151:68:@12512.4]
  assign _T_14730 = entriesToCheck_2_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12514.4]
  assign _T_14731 = _T_14730 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12515.4]
  assign _T_14732 = addrQ_2 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12516.4]
  assign conflict_2_13 = _T_14731 & _T_14732; // @[AxiLoadQueue.scala 151:68:@12517.4]
  assign _T_14734 = entriesToCheck_2_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12519.4]
  assign _T_14735 = _T_14734 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12520.4]
  assign _T_14736 = addrQ_2 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12521.4]
  assign conflict_2_14 = _T_14735 & _T_14736; // @[AxiLoadQueue.scala 151:68:@12522.4]
  assign _T_14738 = entriesToCheck_2_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12524.4]
  assign _T_14739 = _T_14738 & addrKnown_2; // @[AxiLoadQueue.scala 151:41:@12525.4]
  assign _T_14740 = addrQ_2 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12526.4]
  assign conflict_2_15 = _T_14739 & _T_14740; // @[AxiLoadQueue.scala 151:68:@12527.4]
  assign _T_14742 = entriesToCheck_3_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12529.4]
  assign _T_14743 = _T_14742 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12530.4]
  assign _T_14744 = addrQ_3 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12531.4]
  assign conflict_3_0 = _T_14743 & _T_14744; // @[AxiLoadQueue.scala 151:68:@12532.4]
  assign _T_14746 = entriesToCheck_3_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12534.4]
  assign _T_14747 = _T_14746 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12535.4]
  assign _T_14748 = addrQ_3 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12536.4]
  assign conflict_3_1 = _T_14747 & _T_14748; // @[AxiLoadQueue.scala 151:68:@12537.4]
  assign _T_14750 = entriesToCheck_3_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12539.4]
  assign _T_14751 = _T_14750 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12540.4]
  assign _T_14752 = addrQ_3 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12541.4]
  assign conflict_3_2 = _T_14751 & _T_14752; // @[AxiLoadQueue.scala 151:68:@12542.4]
  assign _T_14754 = entriesToCheck_3_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12544.4]
  assign _T_14755 = _T_14754 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12545.4]
  assign _T_14756 = addrQ_3 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12546.4]
  assign conflict_3_3 = _T_14755 & _T_14756; // @[AxiLoadQueue.scala 151:68:@12547.4]
  assign _T_14758 = entriesToCheck_3_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12549.4]
  assign _T_14759 = _T_14758 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12550.4]
  assign _T_14760 = addrQ_3 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12551.4]
  assign conflict_3_4 = _T_14759 & _T_14760; // @[AxiLoadQueue.scala 151:68:@12552.4]
  assign _T_14762 = entriesToCheck_3_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12554.4]
  assign _T_14763 = _T_14762 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12555.4]
  assign _T_14764 = addrQ_3 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12556.4]
  assign conflict_3_5 = _T_14763 & _T_14764; // @[AxiLoadQueue.scala 151:68:@12557.4]
  assign _T_14766 = entriesToCheck_3_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12559.4]
  assign _T_14767 = _T_14766 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12560.4]
  assign _T_14768 = addrQ_3 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12561.4]
  assign conflict_3_6 = _T_14767 & _T_14768; // @[AxiLoadQueue.scala 151:68:@12562.4]
  assign _T_14770 = entriesToCheck_3_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12564.4]
  assign _T_14771 = _T_14770 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12565.4]
  assign _T_14772 = addrQ_3 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12566.4]
  assign conflict_3_7 = _T_14771 & _T_14772; // @[AxiLoadQueue.scala 151:68:@12567.4]
  assign _T_14774 = entriesToCheck_3_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12569.4]
  assign _T_14775 = _T_14774 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12570.4]
  assign _T_14776 = addrQ_3 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12571.4]
  assign conflict_3_8 = _T_14775 & _T_14776; // @[AxiLoadQueue.scala 151:68:@12572.4]
  assign _T_14778 = entriesToCheck_3_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12574.4]
  assign _T_14779 = _T_14778 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12575.4]
  assign _T_14780 = addrQ_3 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12576.4]
  assign conflict_3_9 = _T_14779 & _T_14780; // @[AxiLoadQueue.scala 151:68:@12577.4]
  assign _T_14782 = entriesToCheck_3_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12579.4]
  assign _T_14783 = _T_14782 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12580.4]
  assign _T_14784 = addrQ_3 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12581.4]
  assign conflict_3_10 = _T_14783 & _T_14784; // @[AxiLoadQueue.scala 151:68:@12582.4]
  assign _T_14786 = entriesToCheck_3_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12584.4]
  assign _T_14787 = _T_14786 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12585.4]
  assign _T_14788 = addrQ_3 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12586.4]
  assign conflict_3_11 = _T_14787 & _T_14788; // @[AxiLoadQueue.scala 151:68:@12587.4]
  assign _T_14790 = entriesToCheck_3_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12589.4]
  assign _T_14791 = _T_14790 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12590.4]
  assign _T_14792 = addrQ_3 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12591.4]
  assign conflict_3_12 = _T_14791 & _T_14792; // @[AxiLoadQueue.scala 151:68:@12592.4]
  assign _T_14794 = entriesToCheck_3_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12594.4]
  assign _T_14795 = _T_14794 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12595.4]
  assign _T_14796 = addrQ_3 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12596.4]
  assign conflict_3_13 = _T_14795 & _T_14796; // @[AxiLoadQueue.scala 151:68:@12597.4]
  assign _T_14798 = entriesToCheck_3_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12599.4]
  assign _T_14799 = _T_14798 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12600.4]
  assign _T_14800 = addrQ_3 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12601.4]
  assign conflict_3_14 = _T_14799 & _T_14800; // @[AxiLoadQueue.scala 151:68:@12602.4]
  assign _T_14802 = entriesToCheck_3_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12604.4]
  assign _T_14803 = _T_14802 & addrKnown_3; // @[AxiLoadQueue.scala 151:41:@12605.4]
  assign _T_14804 = addrQ_3 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12606.4]
  assign conflict_3_15 = _T_14803 & _T_14804; // @[AxiLoadQueue.scala 151:68:@12607.4]
  assign _T_14806 = entriesToCheck_4_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12609.4]
  assign _T_14807 = _T_14806 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12610.4]
  assign _T_14808 = addrQ_4 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12611.4]
  assign conflict_4_0 = _T_14807 & _T_14808; // @[AxiLoadQueue.scala 151:68:@12612.4]
  assign _T_14810 = entriesToCheck_4_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12614.4]
  assign _T_14811 = _T_14810 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12615.4]
  assign _T_14812 = addrQ_4 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12616.4]
  assign conflict_4_1 = _T_14811 & _T_14812; // @[AxiLoadQueue.scala 151:68:@12617.4]
  assign _T_14814 = entriesToCheck_4_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12619.4]
  assign _T_14815 = _T_14814 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12620.4]
  assign _T_14816 = addrQ_4 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12621.4]
  assign conflict_4_2 = _T_14815 & _T_14816; // @[AxiLoadQueue.scala 151:68:@12622.4]
  assign _T_14818 = entriesToCheck_4_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12624.4]
  assign _T_14819 = _T_14818 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12625.4]
  assign _T_14820 = addrQ_4 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12626.4]
  assign conflict_4_3 = _T_14819 & _T_14820; // @[AxiLoadQueue.scala 151:68:@12627.4]
  assign _T_14822 = entriesToCheck_4_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12629.4]
  assign _T_14823 = _T_14822 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12630.4]
  assign _T_14824 = addrQ_4 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12631.4]
  assign conflict_4_4 = _T_14823 & _T_14824; // @[AxiLoadQueue.scala 151:68:@12632.4]
  assign _T_14826 = entriesToCheck_4_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12634.4]
  assign _T_14827 = _T_14826 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12635.4]
  assign _T_14828 = addrQ_4 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12636.4]
  assign conflict_4_5 = _T_14827 & _T_14828; // @[AxiLoadQueue.scala 151:68:@12637.4]
  assign _T_14830 = entriesToCheck_4_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12639.4]
  assign _T_14831 = _T_14830 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12640.4]
  assign _T_14832 = addrQ_4 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12641.4]
  assign conflict_4_6 = _T_14831 & _T_14832; // @[AxiLoadQueue.scala 151:68:@12642.4]
  assign _T_14834 = entriesToCheck_4_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12644.4]
  assign _T_14835 = _T_14834 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12645.4]
  assign _T_14836 = addrQ_4 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12646.4]
  assign conflict_4_7 = _T_14835 & _T_14836; // @[AxiLoadQueue.scala 151:68:@12647.4]
  assign _T_14838 = entriesToCheck_4_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12649.4]
  assign _T_14839 = _T_14838 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12650.4]
  assign _T_14840 = addrQ_4 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12651.4]
  assign conflict_4_8 = _T_14839 & _T_14840; // @[AxiLoadQueue.scala 151:68:@12652.4]
  assign _T_14842 = entriesToCheck_4_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12654.4]
  assign _T_14843 = _T_14842 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12655.4]
  assign _T_14844 = addrQ_4 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12656.4]
  assign conflict_4_9 = _T_14843 & _T_14844; // @[AxiLoadQueue.scala 151:68:@12657.4]
  assign _T_14846 = entriesToCheck_4_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12659.4]
  assign _T_14847 = _T_14846 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12660.4]
  assign _T_14848 = addrQ_4 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12661.4]
  assign conflict_4_10 = _T_14847 & _T_14848; // @[AxiLoadQueue.scala 151:68:@12662.4]
  assign _T_14850 = entriesToCheck_4_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12664.4]
  assign _T_14851 = _T_14850 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12665.4]
  assign _T_14852 = addrQ_4 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12666.4]
  assign conflict_4_11 = _T_14851 & _T_14852; // @[AxiLoadQueue.scala 151:68:@12667.4]
  assign _T_14854 = entriesToCheck_4_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12669.4]
  assign _T_14855 = _T_14854 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12670.4]
  assign _T_14856 = addrQ_4 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12671.4]
  assign conflict_4_12 = _T_14855 & _T_14856; // @[AxiLoadQueue.scala 151:68:@12672.4]
  assign _T_14858 = entriesToCheck_4_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12674.4]
  assign _T_14859 = _T_14858 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12675.4]
  assign _T_14860 = addrQ_4 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12676.4]
  assign conflict_4_13 = _T_14859 & _T_14860; // @[AxiLoadQueue.scala 151:68:@12677.4]
  assign _T_14862 = entriesToCheck_4_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12679.4]
  assign _T_14863 = _T_14862 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12680.4]
  assign _T_14864 = addrQ_4 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12681.4]
  assign conflict_4_14 = _T_14863 & _T_14864; // @[AxiLoadQueue.scala 151:68:@12682.4]
  assign _T_14866 = entriesToCheck_4_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12684.4]
  assign _T_14867 = _T_14866 & addrKnown_4; // @[AxiLoadQueue.scala 151:41:@12685.4]
  assign _T_14868 = addrQ_4 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12686.4]
  assign conflict_4_15 = _T_14867 & _T_14868; // @[AxiLoadQueue.scala 151:68:@12687.4]
  assign _T_14870 = entriesToCheck_5_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12689.4]
  assign _T_14871 = _T_14870 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12690.4]
  assign _T_14872 = addrQ_5 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12691.4]
  assign conflict_5_0 = _T_14871 & _T_14872; // @[AxiLoadQueue.scala 151:68:@12692.4]
  assign _T_14874 = entriesToCheck_5_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12694.4]
  assign _T_14875 = _T_14874 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12695.4]
  assign _T_14876 = addrQ_5 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12696.4]
  assign conflict_5_1 = _T_14875 & _T_14876; // @[AxiLoadQueue.scala 151:68:@12697.4]
  assign _T_14878 = entriesToCheck_5_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12699.4]
  assign _T_14879 = _T_14878 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12700.4]
  assign _T_14880 = addrQ_5 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12701.4]
  assign conflict_5_2 = _T_14879 & _T_14880; // @[AxiLoadQueue.scala 151:68:@12702.4]
  assign _T_14882 = entriesToCheck_5_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12704.4]
  assign _T_14883 = _T_14882 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12705.4]
  assign _T_14884 = addrQ_5 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12706.4]
  assign conflict_5_3 = _T_14883 & _T_14884; // @[AxiLoadQueue.scala 151:68:@12707.4]
  assign _T_14886 = entriesToCheck_5_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12709.4]
  assign _T_14887 = _T_14886 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12710.4]
  assign _T_14888 = addrQ_5 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12711.4]
  assign conflict_5_4 = _T_14887 & _T_14888; // @[AxiLoadQueue.scala 151:68:@12712.4]
  assign _T_14890 = entriesToCheck_5_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12714.4]
  assign _T_14891 = _T_14890 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12715.4]
  assign _T_14892 = addrQ_5 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12716.4]
  assign conflict_5_5 = _T_14891 & _T_14892; // @[AxiLoadQueue.scala 151:68:@12717.4]
  assign _T_14894 = entriesToCheck_5_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12719.4]
  assign _T_14895 = _T_14894 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12720.4]
  assign _T_14896 = addrQ_5 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12721.4]
  assign conflict_5_6 = _T_14895 & _T_14896; // @[AxiLoadQueue.scala 151:68:@12722.4]
  assign _T_14898 = entriesToCheck_5_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12724.4]
  assign _T_14899 = _T_14898 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12725.4]
  assign _T_14900 = addrQ_5 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12726.4]
  assign conflict_5_7 = _T_14899 & _T_14900; // @[AxiLoadQueue.scala 151:68:@12727.4]
  assign _T_14902 = entriesToCheck_5_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12729.4]
  assign _T_14903 = _T_14902 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12730.4]
  assign _T_14904 = addrQ_5 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12731.4]
  assign conflict_5_8 = _T_14903 & _T_14904; // @[AxiLoadQueue.scala 151:68:@12732.4]
  assign _T_14906 = entriesToCheck_5_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12734.4]
  assign _T_14907 = _T_14906 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12735.4]
  assign _T_14908 = addrQ_5 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12736.4]
  assign conflict_5_9 = _T_14907 & _T_14908; // @[AxiLoadQueue.scala 151:68:@12737.4]
  assign _T_14910 = entriesToCheck_5_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12739.4]
  assign _T_14911 = _T_14910 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12740.4]
  assign _T_14912 = addrQ_5 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12741.4]
  assign conflict_5_10 = _T_14911 & _T_14912; // @[AxiLoadQueue.scala 151:68:@12742.4]
  assign _T_14914 = entriesToCheck_5_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12744.4]
  assign _T_14915 = _T_14914 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12745.4]
  assign _T_14916 = addrQ_5 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12746.4]
  assign conflict_5_11 = _T_14915 & _T_14916; // @[AxiLoadQueue.scala 151:68:@12747.4]
  assign _T_14918 = entriesToCheck_5_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12749.4]
  assign _T_14919 = _T_14918 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12750.4]
  assign _T_14920 = addrQ_5 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12751.4]
  assign conflict_5_12 = _T_14919 & _T_14920; // @[AxiLoadQueue.scala 151:68:@12752.4]
  assign _T_14922 = entriesToCheck_5_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12754.4]
  assign _T_14923 = _T_14922 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12755.4]
  assign _T_14924 = addrQ_5 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12756.4]
  assign conflict_5_13 = _T_14923 & _T_14924; // @[AxiLoadQueue.scala 151:68:@12757.4]
  assign _T_14926 = entriesToCheck_5_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12759.4]
  assign _T_14927 = _T_14926 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12760.4]
  assign _T_14928 = addrQ_5 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12761.4]
  assign conflict_5_14 = _T_14927 & _T_14928; // @[AxiLoadQueue.scala 151:68:@12762.4]
  assign _T_14930 = entriesToCheck_5_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12764.4]
  assign _T_14931 = _T_14930 & addrKnown_5; // @[AxiLoadQueue.scala 151:41:@12765.4]
  assign _T_14932 = addrQ_5 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12766.4]
  assign conflict_5_15 = _T_14931 & _T_14932; // @[AxiLoadQueue.scala 151:68:@12767.4]
  assign _T_14934 = entriesToCheck_6_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12769.4]
  assign _T_14935 = _T_14934 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12770.4]
  assign _T_14936 = addrQ_6 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12771.4]
  assign conflict_6_0 = _T_14935 & _T_14936; // @[AxiLoadQueue.scala 151:68:@12772.4]
  assign _T_14938 = entriesToCheck_6_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12774.4]
  assign _T_14939 = _T_14938 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12775.4]
  assign _T_14940 = addrQ_6 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12776.4]
  assign conflict_6_1 = _T_14939 & _T_14940; // @[AxiLoadQueue.scala 151:68:@12777.4]
  assign _T_14942 = entriesToCheck_6_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12779.4]
  assign _T_14943 = _T_14942 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12780.4]
  assign _T_14944 = addrQ_6 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12781.4]
  assign conflict_6_2 = _T_14943 & _T_14944; // @[AxiLoadQueue.scala 151:68:@12782.4]
  assign _T_14946 = entriesToCheck_6_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12784.4]
  assign _T_14947 = _T_14946 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12785.4]
  assign _T_14948 = addrQ_6 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12786.4]
  assign conflict_6_3 = _T_14947 & _T_14948; // @[AxiLoadQueue.scala 151:68:@12787.4]
  assign _T_14950 = entriesToCheck_6_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12789.4]
  assign _T_14951 = _T_14950 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12790.4]
  assign _T_14952 = addrQ_6 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12791.4]
  assign conflict_6_4 = _T_14951 & _T_14952; // @[AxiLoadQueue.scala 151:68:@12792.4]
  assign _T_14954 = entriesToCheck_6_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12794.4]
  assign _T_14955 = _T_14954 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12795.4]
  assign _T_14956 = addrQ_6 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12796.4]
  assign conflict_6_5 = _T_14955 & _T_14956; // @[AxiLoadQueue.scala 151:68:@12797.4]
  assign _T_14958 = entriesToCheck_6_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12799.4]
  assign _T_14959 = _T_14958 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12800.4]
  assign _T_14960 = addrQ_6 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12801.4]
  assign conflict_6_6 = _T_14959 & _T_14960; // @[AxiLoadQueue.scala 151:68:@12802.4]
  assign _T_14962 = entriesToCheck_6_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12804.4]
  assign _T_14963 = _T_14962 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12805.4]
  assign _T_14964 = addrQ_6 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12806.4]
  assign conflict_6_7 = _T_14963 & _T_14964; // @[AxiLoadQueue.scala 151:68:@12807.4]
  assign _T_14966 = entriesToCheck_6_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12809.4]
  assign _T_14967 = _T_14966 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12810.4]
  assign _T_14968 = addrQ_6 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12811.4]
  assign conflict_6_8 = _T_14967 & _T_14968; // @[AxiLoadQueue.scala 151:68:@12812.4]
  assign _T_14970 = entriesToCheck_6_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12814.4]
  assign _T_14971 = _T_14970 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12815.4]
  assign _T_14972 = addrQ_6 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12816.4]
  assign conflict_6_9 = _T_14971 & _T_14972; // @[AxiLoadQueue.scala 151:68:@12817.4]
  assign _T_14974 = entriesToCheck_6_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12819.4]
  assign _T_14975 = _T_14974 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12820.4]
  assign _T_14976 = addrQ_6 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12821.4]
  assign conflict_6_10 = _T_14975 & _T_14976; // @[AxiLoadQueue.scala 151:68:@12822.4]
  assign _T_14978 = entriesToCheck_6_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12824.4]
  assign _T_14979 = _T_14978 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12825.4]
  assign _T_14980 = addrQ_6 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12826.4]
  assign conflict_6_11 = _T_14979 & _T_14980; // @[AxiLoadQueue.scala 151:68:@12827.4]
  assign _T_14982 = entriesToCheck_6_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12829.4]
  assign _T_14983 = _T_14982 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12830.4]
  assign _T_14984 = addrQ_6 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12831.4]
  assign conflict_6_12 = _T_14983 & _T_14984; // @[AxiLoadQueue.scala 151:68:@12832.4]
  assign _T_14986 = entriesToCheck_6_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12834.4]
  assign _T_14987 = _T_14986 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12835.4]
  assign _T_14988 = addrQ_6 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12836.4]
  assign conflict_6_13 = _T_14987 & _T_14988; // @[AxiLoadQueue.scala 151:68:@12837.4]
  assign _T_14990 = entriesToCheck_6_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12839.4]
  assign _T_14991 = _T_14990 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12840.4]
  assign _T_14992 = addrQ_6 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12841.4]
  assign conflict_6_14 = _T_14991 & _T_14992; // @[AxiLoadQueue.scala 151:68:@12842.4]
  assign _T_14994 = entriesToCheck_6_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12844.4]
  assign _T_14995 = _T_14994 & addrKnown_6; // @[AxiLoadQueue.scala 151:41:@12845.4]
  assign _T_14996 = addrQ_6 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12846.4]
  assign conflict_6_15 = _T_14995 & _T_14996; // @[AxiLoadQueue.scala 151:68:@12847.4]
  assign _T_14998 = entriesToCheck_7_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12849.4]
  assign _T_14999 = _T_14998 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12850.4]
  assign _T_15000 = addrQ_7 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12851.4]
  assign conflict_7_0 = _T_14999 & _T_15000; // @[AxiLoadQueue.scala 151:68:@12852.4]
  assign _T_15002 = entriesToCheck_7_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12854.4]
  assign _T_15003 = _T_15002 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12855.4]
  assign _T_15004 = addrQ_7 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12856.4]
  assign conflict_7_1 = _T_15003 & _T_15004; // @[AxiLoadQueue.scala 151:68:@12857.4]
  assign _T_15006 = entriesToCheck_7_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12859.4]
  assign _T_15007 = _T_15006 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12860.4]
  assign _T_15008 = addrQ_7 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12861.4]
  assign conflict_7_2 = _T_15007 & _T_15008; // @[AxiLoadQueue.scala 151:68:@12862.4]
  assign _T_15010 = entriesToCheck_7_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12864.4]
  assign _T_15011 = _T_15010 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12865.4]
  assign _T_15012 = addrQ_7 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12866.4]
  assign conflict_7_3 = _T_15011 & _T_15012; // @[AxiLoadQueue.scala 151:68:@12867.4]
  assign _T_15014 = entriesToCheck_7_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12869.4]
  assign _T_15015 = _T_15014 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12870.4]
  assign _T_15016 = addrQ_7 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12871.4]
  assign conflict_7_4 = _T_15015 & _T_15016; // @[AxiLoadQueue.scala 151:68:@12872.4]
  assign _T_15018 = entriesToCheck_7_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12874.4]
  assign _T_15019 = _T_15018 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12875.4]
  assign _T_15020 = addrQ_7 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12876.4]
  assign conflict_7_5 = _T_15019 & _T_15020; // @[AxiLoadQueue.scala 151:68:@12877.4]
  assign _T_15022 = entriesToCheck_7_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12879.4]
  assign _T_15023 = _T_15022 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12880.4]
  assign _T_15024 = addrQ_7 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12881.4]
  assign conflict_7_6 = _T_15023 & _T_15024; // @[AxiLoadQueue.scala 151:68:@12882.4]
  assign _T_15026 = entriesToCheck_7_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12884.4]
  assign _T_15027 = _T_15026 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12885.4]
  assign _T_15028 = addrQ_7 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12886.4]
  assign conflict_7_7 = _T_15027 & _T_15028; // @[AxiLoadQueue.scala 151:68:@12887.4]
  assign _T_15030 = entriesToCheck_7_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12889.4]
  assign _T_15031 = _T_15030 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12890.4]
  assign _T_15032 = addrQ_7 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12891.4]
  assign conflict_7_8 = _T_15031 & _T_15032; // @[AxiLoadQueue.scala 151:68:@12892.4]
  assign _T_15034 = entriesToCheck_7_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12894.4]
  assign _T_15035 = _T_15034 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12895.4]
  assign _T_15036 = addrQ_7 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12896.4]
  assign conflict_7_9 = _T_15035 & _T_15036; // @[AxiLoadQueue.scala 151:68:@12897.4]
  assign _T_15038 = entriesToCheck_7_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12899.4]
  assign _T_15039 = _T_15038 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12900.4]
  assign _T_15040 = addrQ_7 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12901.4]
  assign conflict_7_10 = _T_15039 & _T_15040; // @[AxiLoadQueue.scala 151:68:@12902.4]
  assign _T_15042 = entriesToCheck_7_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12904.4]
  assign _T_15043 = _T_15042 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12905.4]
  assign _T_15044 = addrQ_7 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12906.4]
  assign conflict_7_11 = _T_15043 & _T_15044; // @[AxiLoadQueue.scala 151:68:@12907.4]
  assign _T_15046 = entriesToCheck_7_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12909.4]
  assign _T_15047 = _T_15046 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12910.4]
  assign _T_15048 = addrQ_7 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12911.4]
  assign conflict_7_12 = _T_15047 & _T_15048; // @[AxiLoadQueue.scala 151:68:@12912.4]
  assign _T_15050 = entriesToCheck_7_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12914.4]
  assign _T_15051 = _T_15050 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12915.4]
  assign _T_15052 = addrQ_7 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12916.4]
  assign conflict_7_13 = _T_15051 & _T_15052; // @[AxiLoadQueue.scala 151:68:@12917.4]
  assign _T_15054 = entriesToCheck_7_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12919.4]
  assign _T_15055 = _T_15054 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12920.4]
  assign _T_15056 = addrQ_7 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@12921.4]
  assign conflict_7_14 = _T_15055 & _T_15056; // @[AxiLoadQueue.scala 151:68:@12922.4]
  assign _T_15058 = entriesToCheck_7_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@12924.4]
  assign _T_15059 = _T_15058 & addrKnown_7; // @[AxiLoadQueue.scala 151:41:@12925.4]
  assign _T_15060 = addrQ_7 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@12926.4]
  assign conflict_7_15 = _T_15059 & _T_15060; // @[AxiLoadQueue.scala 151:68:@12927.4]
  assign _T_15062 = entriesToCheck_8_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@12929.4]
  assign _T_15063 = _T_15062 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12930.4]
  assign _T_15064 = addrQ_8 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@12931.4]
  assign conflict_8_0 = _T_15063 & _T_15064; // @[AxiLoadQueue.scala 151:68:@12932.4]
  assign _T_15066 = entriesToCheck_8_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@12934.4]
  assign _T_15067 = _T_15066 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12935.4]
  assign _T_15068 = addrQ_8 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@12936.4]
  assign conflict_8_1 = _T_15067 & _T_15068; // @[AxiLoadQueue.scala 151:68:@12937.4]
  assign _T_15070 = entriesToCheck_8_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@12939.4]
  assign _T_15071 = _T_15070 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12940.4]
  assign _T_15072 = addrQ_8 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@12941.4]
  assign conflict_8_2 = _T_15071 & _T_15072; // @[AxiLoadQueue.scala 151:68:@12942.4]
  assign _T_15074 = entriesToCheck_8_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@12944.4]
  assign _T_15075 = _T_15074 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12945.4]
  assign _T_15076 = addrQ_8 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@12946.4]
  assign conflict_8_3 = _T_15075 & _T_15076; // @[AxiLoadQueue.scala 151:68:@12947.4]
  assign _T_15078 = entriesToCheck_8_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@12949.4]
  assign _T_15079 = _T_15078 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12950.4]
  assign _T_15080 = addrQ_8 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@12951.4]
  assign conflict_8_4 = _T_15079 & _T_15080; // @[AxiLoadQueue.scala 151:68:@12952.4]
  assign _T_15082 = entriesToCheck_8_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@12954.4]
  assign _T_15083 = _T_15082 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12955.4]
  assign _T_15084 = addrQ_8 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@12956.4]
  assign conflict_8_5 = _T_15083 & _T_15084; // @[AxiLoadQueue.scala 151:68:@12957.4]
  assign _T_15086 = entriesToCheck_8_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@12959.4]
  assign _T_15087 = _T_15086 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12960.4]
  assign _T_15088 = addrQ_8 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@12961.4]
  assign conflict_8_6 = _T_15087 & _T_15088; // @[AxiLoadQueue.scala 151:68:@12962.4]
  assign _T_15090 = entriesToCheck_8_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@12964.4]
  assign _T_15091 = _T_15090 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12965.4]
  assign _T_15092 = addrQ_8 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@12966.4]
  assign conflict_8_7 = _T_15091 & _T_15092; // @[AxiLoadQueue.scala 151:68:@12967.4]
  assign _T_15094 = entriesToCheck_8_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@12969.4]
  assign _T_15095 = _T_15094 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12970.4]
  assign _T_15096 = addrQ_8 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@12971.4]
  assign conflict_8_8 = _T_15095 & _T_15096; // @[AxiLoadQueue.scala 151:68:@12972.4]
  assign _T_15098 = entriesToCheck_8_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@12974.4]
  assign _T_15099 = _T_15098 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12975.4]
  assign _T_15100 = addrQ_8 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@12976.4]
  assign conflict_8_9 = _T_15099 & _T_15100; // @[AxiLoadQueue.scala 151:68:@12977.4]
  assign _T_15102 = entriesToCheck_8_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@12979.4]
  assign _T_15103 = _T_15102 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12980.4]
  assign _T_15104 = addrQ_8 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@12981.4]
  assign conflict_8_10 = _T_15103 & _T_15104; // @[AxiLoadQueue.scala 151:68:@12982.4]
  assign _T_15106 = entriesToCheck_8_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@12984.4]
  assign _T_15107 = _T_15106 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12985.4]
  assign _T_15108 = addrQ_8 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@12986.4]
  assign conflict_8_11 = _T_15107 & _T_15108; // @[AxiLoadQueue.scala 151:68:@12987.4]
  assign _T_15110 = entriesToCheck_8_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@12989.4]
  assign _T_15111 = _T_15110 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12990.4]
  assign _T_15112 = addrQ_8 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@12991.4]
  assign conflict_8_12 = _T_15111 & _T_15112; // @[AxiLoadQueue.scala 151:68:@12992.4]
  assign _T_15114 = entriesToCheck_8_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@12994.4]
  assign _T_15115 = _T_15114 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@12995.4]
  assign _T_15116 = addrQ_8 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@12996.4]
  assign conflict_8_13 = _T_15115 & _T_15116; // @[AxiLoadQueue.scala 151:68:@12997.4]
  assign _T_15118 = entriesToCheck_8_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@12999.4]
  assign _T_15119 = _T_15118 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@13000.4]
  assign _T_15120 = addrQ_8 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13001.4]
  assign conflict_8_14 = _T_15119 & _T_15120; // @[AxiLoadQueue.scala 151:68:@13002.4]
  assign _T_15122 = entriesToCheck_8_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13004.4]
  assign _T_15123 = _T_15122 & addrKnown_8; // @[AxiLoadQueue.scala 151:41:@13005.4]
  assign _T_15124 = addrQ_8 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13006.4]
  assign conflict_8_15 = _T_15123 & _T_15124; // @[AxiLoadQueue.scala 151:68:@13007.4]
  assign _T_15126 = entriesToCheck_9_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@13009.4]
  assign _T_15127 = _T_15126 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13010.4]
  assign _T_15128 = addrQ_9 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@13011.4]
  assign conflict_9_0 = _T_15127 & _T_15128; // @[AxiLoadQueue.scala 151:68:@13012.4]
  assign _T_15130 = entriesToCheck_9_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@13014.4]
  assign _T_15131 = _T_15130 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13015.4]
  assign _T_15132 = addrQ_9 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@13016.4]
  assign conflict_9_1 = _T_15131 & _T_15132; // @[AxiLoadQueue.scala 151:68:@13017.4]
  assign _T_15134 = entriesToCheck_9_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@13019.4]
  assign _T_15135 = _T_15134 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13020.4]
  assign _T_15136 = addrQ_9 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@13021.4]
  assign conflict_9_2 = _T_15135 & _T_15136; // @[AxiLoadQueue.scala 151:68:@13022.4]
  assign _T_15138 = entriesToCheck_9_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@13024.4]
  assign _T_15139 = _T_15138 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13025.4]
  assign _T_15140 = addrQ_9 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@13026.4]
  assign conflict_9_3 = _T_15139 & _T_15140; // @[AxiLoadQueue.scala 151:68:@13027.4]
  assign _T_15142 = entriesToCheck_9_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@13029.4]
  assign _T_15143 = _T_15142 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13030.4]
  assign _T_15144 = addrQ_9 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@13031.4]
  assign conflict_9_4 = _T_15143 & _T_15144; // @[AxiLoadQueue.scala 151:68:@13032.4]
  assign _T_15146 = entriesToCheck_9_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@13034.4]
  assign _T_15147 = _T_15146 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13035.4]
  assign _T_15148 = addrQ_9 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@13036.4]
  assign conflict_9_5 = _T_15147 & _T_15148; // @[AxiLoadQueue.scala 151:68:@13037.4]
  assign _T_15150 = entriesToCheck_9_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@13039.4]
  assign _T_15151 = _T_15150 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13040.4]
  assign _T_15152 = addrQ_9 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@13041.4]
  assign conflict_9_6 = _T_15151 & _T_15152; // @[AxiLoadQueue.scala 151:68:@13042.4]
  assign _T_15154 = entriesToCheck_9_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@13044.4]
  assign _T_15155 = _T_15154 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13045.4]
  assign _T_15156 = addrQ_9 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@13046.4]
  assign conflict_9_7 = _T_15155 & _T_15156; // @[AxiLoadQueue.scala 151:68:@13047.4]
  assign _T_15158 = entriesToCheck_9_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@13049.4]
  assign _T_15159 = _T_15158 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13050.4]
  assign _T_15160 = addrQ_9 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@13051.4]
  assign conflict_9_8 = _T_15159 & _T_15160; // @[AxiLoadQueue.scala 151:68:@13052.4]
  assign _T_15162 = entriesToCheck_9_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@13054.4]
  assign _T_15163 = _T_15162 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13055.4]
  assign _T_15164 = addrQ_9 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@13056.4]
  assign conflict_9_9 = _T_15163 & _T_15164; // @[AxiLoadQueue.scala 151:68:@13057.4]
  assign _T_15166 = entriesToCheck_9_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@13059.4]
  assign _T_15167 = _T_15166 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13060.4]
  assign _T_15168 = addrQ_9 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@13061.4]
  assign conflict_9_10 = _T_15167 & _T_15168; // @[AxiLoadQueue.scala 151:68:@13062.4]
  assign _T_15170 = entriesToCheck_9_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@13064.4]
  assign _T_15171 = _T_15170 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13065.4]
  assign _T_15172 = addrQ_9 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@13066.4]
  assign conflict_9_11 = _T_15171 & _T_15172; // @[AxiLoadQueue.scala 151:68:@13067.4]
  assign _T_15174 = entriesToCheck_9_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@13069.4]
  assign _T_15175 = _T_15174 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13070.4]
  assign _T_15176 = addrQ_9 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@13071.4]
  assign conflict_9_12 = _T_15175 & _T_15176; // @[AxiLoadQueue.scala 151:68:@13072.4]
  assign _T_15178 = entriesToCheck_9_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@13074.4]
  assign _T_15179 = _T_15178 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13075.4]
  assign _T_15180 = addrQ_9 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@13076.4]
  assign conflict_9_13 = _T_15179 & _T_15180; // @[AxiLoadQueue.scala 151:68:@13077.4]
  assign _T_15182 = entriesToCheck_9_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@13079.4]
  assign _T_15183 = _T_15182 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13080.4]
  assign _T_15184 = addrQ_9 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13081.4]
  assign conflict_9_14 = _T_15183 & _T_15184; // @[AxiLoadQueue.scala 151:68:@13082.4]
  assign _T_15186 = entriesToCheck_9_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13084.4]
  assign _T_15187 = _T_15186 & addrKnown_9; // @[AxiLoadQueue.scala 151:41:@13085.4]
  assign _T_15188 = addrQ_9 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13086.4]
  assign conflict_9_15 = _T_15187 & _T_15188; // @[AxiLoadQueue.scala 151:68:@13087.4]
  assign _T_15190 = entriesToCheck_10_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@13089.4]
  assign _T_15191 = _T_15190 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13090.4]
  assign _T_15192 = addrQ_10 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@13091.4]
  assign conflict_10_0 = _T_15191 & _T_15192; // @[AxiLoadQueue.scala 151:68:@13092.4]
  assign _T_15194 = entriesToCheck_10_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@13094.4]
  assign _T_15195 = _T_15194 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13095.4]
  assign _T_15196 = addrQ_10 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@13096.4]
  assign conflict_10_1 = _T_15195 & _T_15196; // @[AxiLoadQueue.scala 151:68:@13097.4]
  assign _T_15198 = entriesToCheck_10_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@13099.4]
  assign _T_15199 = _T_15198 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13100.4]
  assign _T_15200 = addrQ_10 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@13101.4]
  assign conflict_10_2 = _T_15199 & _T_15200; // @[AxiLoadQueue.scala 151:68:@13102.4]
  assign _T_15202 = entriesToCheck_10_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@13104.4]
  assign _T_15203 = _T_15202 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13105.4]
  assign _T_15204 = addrQ_10 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@13106.4]
  assign conflict_10_3 = _T_15203 & _T_15204; // @[AxiLoadQueue.scala 151:68:@13107.4]
  assign _T_15206 = entriesToCheck_10_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@13109.4]
  assign _T_15207 = _T_15206 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13110.4]
  assign _T_15208 = addrQ_10 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@13111.4]
  assign conflict_10_4 = _T_15207 & _T_15208; // @[AxiLoadQueue.scala 151:68:@13112.4]
  assign _T_15210 = entriesToCheck_10_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@13114.4]
  assign _T_15211 = _T_15210 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13115.4]
  assign _T_15212 = addrQ_10 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@13116.4]
  assign conflict_10_5 = _T_15211 & _T_15212; // @[AxiLoadQueue.scala 151:68:@13117.4]
  assign _T_15214 = entriesToCheck_10_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@13119.4]
  assign _T_15215 = _T_15214 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13120.4]
  assign _T_15216 = addrQ_10 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@13121.4]
  assign conflict_10_6 = _T_15215 & _T_15216; // @[AxiLoadQueue.scala 151:68:@13122.4]
  assign _T_15218 = entriesToCheck_10_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@13124.4]
  assign _T_15219 = _T_15218 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13125.4]
  assign _T_15220 = addrQ_10 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@13126.4]
  assign conflict_10_7 = _T_15219 & _T_15220; // @[AxiLoadQueue.scala 151:68:@13127.4]
  assign _T_15222 = entriesToCheck_10_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@13129.4]
  assign _T_15223 = _T_15222 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13130.4]
  assign _T_15224 = addrQ_10 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@13131.4]
  assign conflict_10_8 = _T_15223 & _T_15224; // @[AxiLoadQueue.scala 151:68:@13132.4]
  assign _T_15226 = entriesToCheck_10_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@13134.4]
  assign _T_15227 = _T_15226 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13135.4]
  assign _T_15228 = addrQ_10 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@13136.4]
  assign conflict_10_9 = _T_15227 & _T_15228; // @[AxiLoadQueue.scala 151:68:@13137.4]
  assign _T_15230 = entriesToCheck_10_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@13139.4]
  assign _T_15231 = _T_15230 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13140.4]
  assign _T_15232 = addrQ_10 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@13141.4]
  assign conflict_10_10 = _T_15231 & _T_15232; // @[AxiLoadQueue.scala 151:68:@13142.4]
  assign _T_15234 = entriesToCheck_10_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@13144.4]
  assign _T_15235 = _T_15234 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13145.4]
  assign _T_15236 = addrQ_10 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@13146.4]
  assign conflict_10_11 = _T_15235 & _T_15236; // @[AxiLoadQueue.scala 151:68:@13147.4]
  assign _T_15238 = entriesToCheck_10_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@13149.4]
  assign _T_15239 = _T_15238 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13150.4]
  assign _T_15240 = addrQ_10 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@13151.4]
  assign conflict_10_12 = _T_15239 & _T_15240; // @[AxiLoadQueue.scala 151:68:@13152.4]
  assign _T_15242 = entriesToCheck_10_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@13154.4]
  assign _T_15243 = _T_15242 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13155.4]
  assign _T_15244 = addrQ_10 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@13156.4]
  assign conflict_10_13 = _T_15243 & _T_15244; // @[AxiLoadQueue.scala 151:68:@13157.4]
  assign _T_15246 = entriesToCheck_10_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@13159.4]
  assign _T_15247 = _T_15246 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13160.4]
  assign _T_15248 = addrQ_10 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13161.4]
  assign conflict_10_14 = _T_15247 & _T_15248; // @[AxiLoadQueue.scala 151:68:@13162.4]
  assign _T_15250 = entriesToCheck_10_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13164.4]
  assign _T_15251 = _T_15250 & addrKnown_10; // @[AxiLoadQueue.scala 151:41:@13165.4]
  assign _T_15252 = addrQ_10 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13166.4]
  assign conflict_10_15 = _T_15251 & _T_15252; // @[AxiLoadQueue.scala 151:68:@13167.4]
  assign _T_15254 = entriesToCheck_11_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@13169.4]
  assign _T_15255 = _T_15254 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13170.4]
  assign _T_15256 = addrQ_11 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@13171.4]
  assign conflict_11_0 = _T_15255 & _T_15256; // @[AxiLoadQueue.scala 151:68:@13172.4]
  assign _T_15258 = entriesToCheck_11_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@13174.4]
  assign _T_15259 = _T_15258 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13175.4]
  assign _T_15260 = addrQ_11 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@13176.4]
  assign conflict_11_1 = _T_15259 & _T_15260; // @[AxiLoadQueue.scala 151:68:@13177.4]
  assign _T_15262 = entriesToCheck_11_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@13179.4]
  assign _T_15263 = _T_15262 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13180.4]
  assign _T_15264 = addrQ_11 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@13181.4]
  assign conflict_11_2 = _T_15263 & _T_15264; // @[AxiLoadQueue.scala 151:68:@13182.4]
  assign _T_15266 = entriesToCheck_11_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@13184.4]
  assign _T_15267 = _T_15266 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13185.4]
  assign _T_15268 = addrQ_11 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@13186.4]
  assign conflict_11_3 = _T_15267 & _T_15268; // @[AxiLoadQueue.scala 151:68:@13187.4]
  assign _T_15270 = entriesToCheck_11_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@13189.4]
  assign _T_15271 = _T_15270 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13190.4]
  assign _T_15272 = addrQ_11 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@13191.4]
  assign conflict_11_4 = _T_15271 & _T_15272; // @[AxiLoadQueue.scala 151:68:@13192.4]
  assign _T_15274 = entriesToCheck_11_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@13194.4]
  assign _T_15275 = _T_15274 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13195.4]
  assign _T_15276 = addrQ_11 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@13196.4]
  assign conflict_11_5 = _T_15275 & _T_15276; // @[AxiLoadQueue.scala 151:68:@13197.4]
  assign _T_15278 = entriesToCheck_11_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@13199.4]
  assign _T_15279 = _T_15278 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13200.4]
  assign _T_15280 = addrQ_11 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@13201.4]
  assign conflict_11_6 = _T_15279 & _T_15280; // @[AxiLoadQueue.scala 151:68:@13202.4]
  assign _T_15282 = entriesToCheck_11_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@13204.4]
  assign _T_15283 = _T_15282 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13205.4]
  assign _T_15284 = addrQ_11 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@13206.4]
  assign conflict_11_7 = _T_15283 & _T_15284; // @[AxiLoadQueue.scala 151:68:@13207.4]
  assign _T_15286 = entriesToCheck_11_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@13209.4]
  assign _T_15287 = _T_15286 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13210.4]
  assign _T_15288 = addrQ_11 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@13211.4]
  assign conflict_11_8 = _T_15287 & _T_15288; // @[AxiLoadQueue.scala 151:68:@13212.4]
  assign _T_15290 = entriesToCheck_11_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@13214.4]
  assign _T_15291 = _T_15290 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13215.4]
  assign _T_15292 = addrQ_11 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@13216.4]
  assign conflict_11_9 = _T_15291 & _T_15292; // @[AxiLoadQueue.scala 151:68:@13217.4]
  assign _T_15294 = entriesToCheck_11_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@13219.4]
  assign _T_15295 = _T_15294 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13220.4]
  assign _T_15296 = addrQ_11 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@13221.4]
  assign conflict_11_10 = _T_15295 & _T_15296; // @[AxiLoadQueue.scala 151:68:@13222.4]
  assign _T_15298 = entriesToCheck_11_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@13224.4]
  assign _T_15299 = _T_15298 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13225.4]
  assign _T_15300 = addrQ_11 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@13226.4]
  assign conflict_11_11 = _T_15299 & _T_15300; // @[AxiLoadQueue.scala 151:68:@13227.4]
  assign _T_15302 = entriesToCheck_11_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@13229.4]
  assign _T_15303 = _T_15302 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13230.4]
  assign _T_15304 = addrQ_11 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@13231.4]
  assign conflict_11_12 = _T_15303 & _T_15304; // @[AxiLoadQueue.scala 151:68:@13232.4]
  assign _T_15306 = entriesToCheck_11_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@13234.4]
  assign _T_15307 = _T_15306 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13235.4]
  assign _T_15308 = addrQ_11 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@13236.4]
  assign conflict_11_13 = _T_15307 & _T_15308; // @[AxiLoadQueue.scala 151:68:@13237.4]
  assign _T_15310 = entriesToCheck_11_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@13239.4]
  assign _T_15311 = _T_15310 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13240.4]
  assign _T_15312 = addrQ_11 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13241.4]
  assign conflict_11_14 = _T_15311 & _T_15312; // @[AxiLoadQueue.scala 151:68:@13242.4]
  assign _T_15314 = entriesToCheck_11_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13244.4]
  assign _T_15315 = _T_15314 & addrKnown_11; // @[AxiLoadQueue.scala 151:41:@13245.4]
  assign _T_15316 = addrQ_11 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13246.4]
  assign conflict_11_15 = _T_15315 & _T_15316; // @[AxiLoadQueue.scala 151:68:@13247.4]
  assign _T_15318 = entriesToCheck_12_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@13249.4]
  assign _T_15319 = _T_15318 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13250.4]
  assign _T_15320 = addrQ_12 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@13251.4]
  assign conflict_12_0 = _T_15319 & _T_15320; // @[AxiLoadQueue.scala 151:68:@13252.4]
  assign _T_15322 = entriesToCheck_12_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@13254.4]
  assign _T_15323 = _T_15322 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13255.4]
  assign _T_15324 = addrQ_12 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@13256.4]
  assign conflict_12_1 = _T_15323 & _T_15324; // @[AxiLoadQueue.scala 151:68:@13257.4]
  assign _T_15326 = entriesToCheck_12_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@13259.4]
  assign _T_15327 = _T_15326 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13260.4]
  assign _T_15328 = addrQ_12 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@13261.4]
  assign conflict_12_2 = _T_15327 & _T_15328; // @[AxiLoadQueue.scala 151:68:@13262.4]
  assign _T_15330 = entriesToCheck_12_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@13264.4]
  assign _T_15331 = _T_15330 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13265.4]
  assign _T_15332 = addrQ_12 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@13266.4]
  assign conflict_12_3 = _T_15331 & _T_15332; // @[AxiLoadQueue.scala 151:68:@13267.4]
  assign _T_15334 = entriesToCheck_12_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@13269.4]
  assign _T_15335 = _T_15334 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13270.4]
  assign _T_15336 = addrQ_12 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@13271.4]
  assign conflict_12_4 = _T_15335 & _T_15336; // @[AxiLoadQueue.scala 151:68:@13272.4]
  assign _T_15338 = entriesToCheck_12_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@13274.4]
  assign _T_15339 = _T_15338 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13275.4]
  assign _T_15340 = addrQ_12 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@13276.4]
  assign conflict_12_5 = _T_15339 & _T_15340; // @[AxiLoadQueue.scala 151:68:@13277.4]
  assign _T_15342 = entriesToCheck_12_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@13279.4]
  assign _T_15343 = _T_15342 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13280.4]
  assign _T_15344 = addrQ_12 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@13281.4]
  assign conflict_12_6 = _T_15343 & _T_15344; // @[AxiLoadQueue.scala 151:68:@13282.4]
  assign _T_15346 = entriesToCheck_12_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@13284.4]
  assign _T_15347 = _T_15346 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13285.4]
  assign _T_15348 = addrQ_12 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@13286.4]
  assign conflict_12_7 = _T_15347 & _T_15348; // @[AxiLoadQueue.scala 151:68:@13287.4]
  assign _T_15350 = entriesToCheck_12_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@13289.4]
  assign _T_15351 = _T_15350 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13290.4]
  assign _T_15352 = addrQ_12 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@13291.4]
  assign conflict_12_8 = _T_15351 & _T_15352; // @[AxiLoadQueue.scala 151:68:@13292.4]
  assign _T_15354 = entriesToCheck_12_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@13294.4]
  assign _T_15355 = _T_15354 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13295.4]
  assign _T_15356 = addrQ_12 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@13296.4]
  assign conflict_12_9 = _T_15355 & _T_15356; // @[AxiLoadQueue.scala 151:68:@13297.4]
  assign _T_15358 = entriesToCheck_12_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@13299.4]
  assign _T_15359 = _T_15358 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13300.4]
  assign _T_15360 = addrQ_12 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@13301.4]
  assign conflict_12_10 = _T_15359 & _T_15360; // @[AxiLoadQueue.scala 151:68:@13302.4]
  assign _T_15362 = entriesToCheck_12_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@13304.4]
  assign _T_15363 = _T_15362 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13305.4]
  assign _T_15364 = addrQ_12 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@13306.4]
  assign conflict_12_11 = _T_15363 & _T_15364; // @[AxiLoadQueue.scala 151:68:@13307.4]
  assign _T_15366 = entriesToCheck_12_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@13309.4]
  assign _T_15367 = _T_15366 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13310.4]
  assign _T_15368 = addrQ_12 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@13311.4]
  assign conflict_12_12 = _T_15367 & _T_15368; // @[AxiLoadQueue.scala 151:68:@13312.4]
  assign _T_15370 = entriesToCheck_12_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@13314.4]
  assign _T_15371 = _T_15370 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13315.4]
  assign _T_15372 = addrQ_12 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@13316.4]
  assign conflict_12_13 = _T_15371 & _T_15372; // @[AxiLoadQueue.scala 151:68:@13317.4]
  assign _T_15374 = entriesToCheck_12_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@13319.4]
  assign _T_15375 = _T_15374 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13320.4]
  assign _T_15376 = addrQ_12 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13321.4]
  assign conflict_12_14 = _T_15375 & _T_15376; // @[AxiLoadQueue.scala 151:68:@13322.4]
  assign _T_15378 = entriesToCheck_12_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13324.4]
  assign _T_15379 = _T_15378 & addrKnown_12; // @[AxiLoadQueue.scala 151:41:@13325.4]
  assign _T_15380 = addrQ_12 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13326.4]
  assign conflict_12_15 = _T_15379 & _T_15380; // @[AxiLoadQueue.scala 151:68:@13327.4]
  assign _T_15382 = entriesToCheck_13_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@13329.4]
  assign _T_15383 = _T_15382 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13330.4]
  assign _T_15384 = addrQ_13 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@13331.4]
  assign conflict_13_0 = _T_15383 & _T_15384; // @[AxiLoadQueue.scala 151:68:@13332.4]
  assign _T_15386 = entriesToCheck_13_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@13334.4]
  assign _T_15387 = _T_15386 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13335.4]
  assign _T_15388 = addrQ_13 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@13336.4]
  assign conflict_13_1 = _T_15387 & _T_15388; // @[AxiLoadQueue.scala 151:68:@13337.4]
  assign _T_15390 = entriesToCheck_13_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@13339.4]
  assign _T_15391 = _T_15390 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13340.4]
  assign _T_15392 = addrQ_13 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@13341.4]
  assign conflict_13_2 = _T_15391 & _T_15392; // @[AxiLoadQueue.scala 151:68:@13342.4]
  assign _T_15394 = entriesToCheck_13_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@13344.4]
  assign _T_15395 = _T_15394 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13345.4]
  assign _T_15396 = addrQ_13 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@13346.4]
  assign conflict_13_3 = _T_15395 & _T_15396; // @[AxiLoadQueue.scala 151:68:@13347.4]
  assign _T_15398 = entriesToCheck_13_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@13349.4]
  assign _T_15399 = _T_15398 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13350.4]
  assign _T_15400 = addrQ_13 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@13351.4]
  assign conflict_13_4 = _T_15399 & _T_15400; // @[AxiLoadQueue.scala 151:68:@13352.4]
  assign _T_15402 = entriesToCheck_13_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@13354.4]
  assign _T_15403 = _T_15402 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13355.4]
  assign _T_15404 = addrQ_13 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@13356.4]
  assign conflict_13_5 = _T_15403 & _T_15404; // @[AxiLoadQueue.scala 151:68:@13357.4]
  assign _T_15406 = entriesToCheck_13_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@13359.4]
  assign _T_15407 = _T_15406 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13360.4]
  assign _T_15408 = addrQ_13 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@13361.4]
  assign conflict_13_6 = _T_15407 & _T_15408; // @[AxiLoadQueue.scala 151:68:@13362.4]
  assign _T_15410 = entriesToCheck_13_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@13364.4]
  assign _T_15411 = _T_15410 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13365.4]
  assign _T_15412 = addrQ_13 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@13366.4]
  assign conflict_13_7 = _T_15411 & _T_15412; // @[AxiLoadQueue.scala 151:68:@13367.4]
  assign _T_15414 = entriesToCheck_13_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@13369.4]
  assign _T_15415 = _T_15414 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13370.4]
  assign _T_15416 = addrQ_13 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@13371.4]
  assign conflict_13_8 = _T_15415 & _T_15416; // @[AxiLoadQueue.scala 151:68:@13372.4]
  assign _T_15418 = entriesToCheck_13_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@13374.4]
  assign _T_15419 = _T_15418 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13375.4]
  assign _T_15420 = addrQ_13 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@13376.4]
  assign conflict_13_9 = _T_15419 & _T_15420; // @[AxiLoadQueue.scala 151:68:@13377.4]
  assign _T_15422 = entriesToCheck_13_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@13379.4]
  assign _T_15423 = _T_15422 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13380.4]
  assign _T_15424 = addrQ_13 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@13381.4]
  assign conflict_13_10 = _T_15423 & _T_15424; // @[AxiLoadQueue.scala 151:68:@13382.4]
  assign _T_15426 = entriesToCheck_13_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@13384.4]
  assign _T_15427 = _T_15426 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13385.4]
  assign _T_15428 = addrQ_13 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@13386.4]
  assign conflict_13_11 = _T_15427 & _T_15428; // @[AxiLoadQueue.scala 151:68:@13387.4]
  assign _T_15430 = entriesToCheck_13_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@13389.4]
  assign _T_15431 = _T_15430 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13390.4]
  assign _T_15432 = addrQ_13 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@13391.4]
  assign conflict_13_12 = _T_15431 & _T_15432; // @[AxiLoadQueue.scala 151:68:@13392.4]
  assign _T_15434 = entriesToCheck_13_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@13394.4]
  assign _T_15435 = _T_15434 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13395.4]
  assign _T_15436 = addrQ_13 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@13396.4]
  assign conflict_13_13 = _T_15435 & _T_15436; // @[AxiLoadQueue.scala 151:68:@13397.4]
  assign _T_15438 = entriesToCheck_13_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@13399.4]
  assign _T_15439 = _T_15438 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13400.4]
  assign _T_15440 = addrQ_13 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13401.4]
  assign conflict_13_14 = _T_15439 & _T_15440; // @[AxiLoadQueue.scala 151:68:@13402.4]
  assign _T_15442 = entriesToCheck_13_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13404.4]
  assign _T_15443 = _T_15442 & addrKnown_13; // @[AxiLoadQueue.scala 151:41:@13405.4]
  assign _T_15444 = addrQ_13 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13406.4]
  assign conflict_13_15 = _T_15443 & _T_15444; // @[AxiLoadQueue.scala 151:68:@13407.4]
  assign _T_15446 = entriesToCheck_14_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@13409.4]
  assign _T_15447 = _T_15446 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13410.4]
  assign _T_15448 = addrQ_14 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@13411.4]
  assign conflict_14_0 = _T_15447 & _T_15448; // @[AxiLoadQueue.scala 151:68:@13412.4]
  assign _T_15450 = entriesToCheck_14_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@13414.4]
  assign _T_15451 = _T_15450 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13415.4]
  assign _T_15452 = addrQ_14 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@13416.4]
  assign conflict_14_1 = _T_15451 & _T_15452; // @[AxiLoadQueue.scala 151:68:@13417.4]
  assign _T_15454 = entriesToCheck_14_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@13419.4]
  assign _T_15455 = _T_15454 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13420.4]
  assign _T_15456 = addrQ_14 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@13421.4]
  assign conflict_14_2 = _T_15455 & _T_15456; // @[AxiLoadQueue.scala 151:68:@13422.4]
  assign _T_15458 = entriesToCheck_14_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@13424.4]
  assign _T_15459 = _T_15458 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13425.4]
  assign _T_15460 = addrQ_14 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@13426.4]
  assign conflict_14_3 = _T_15459 & _T_15460; // @[AxiLoadQueue.scala 151:68:@13427.4]
  assign _T_15462 = entriesToCheck_14_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@13429.4]
  assign _T_15463 = _T_15462 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13430.4]
  assign _T_15464 = addrQ_14 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@13431.4]
  assign conflict_14_4 = _T_15463 & _T_15464; // @[AxiLoadQueue.scala 151:68:@13432.4]
  assign _T_15466 = entriesToCheck_14_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@13434.4]
  assign _T_15467 = _T_15466 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13435.4]
  assign _T_15468 = addrQ_14 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@13436.4]
  assign conflict_14_5 = _T_15467 & _T_15468; // @[AxiLoadQueue.scala 151:68:@13437.4]
  assign _T_15470 = entriesToCheck_14_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@13439.4]
  assign _T_15471 = _T_15470 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13440.4]
  assign _T_15472 = addrQ_14 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@13441.4]
  assign conflict_14_6 = _T_15471 & _T_15472; // @[AxiLoadQueue.scala 151:68:@13442.4]
  assign _T_15474 = entriesToCheck_14_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@13444.4]
  assign _T_15475 = _T_15474 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13445.4]
  assign _T_15476 = addrQ_14 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@13446.4]
  assign conflict_14_7 = _T_15475 & _T_15476; // @[AxiLoadQueue.scala 151:68:@13447.4]
  assign _T_15478 = entriesToCheck_14_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@13449.4]
  assign _T_15479 = _T_15478 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13450.4]
  assign _T_15480 = addrQ_14 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@13451.4]
  assign conflict_14_8 = _T_15479 & _T_15480; // @[AxiLoadQueue.scala 151:68:@13452.4]
  assign _T_15482 = entriesToCheck_14_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@13454.4]
  assign _T_15483 = _T_15482 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13455.4]
  assign _T_15484 = addrQ_14 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@13456.4]
  assign conflict_14_9 = _T_15483 & _T_15484; // @[AxiLoadQueue.scala 151:68:@13457.4]
  assign _T_15486 = entriesToCheck_14_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@13459.4]
  assign _T_15487 = _T_15486 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13460.4]
  assign _T_15488 = addrQ_14 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@13461.4]
  assign conflict_14_10 = _T_15487 & _T_15488; // @[AxiLoadQueue.scala 151:68:@13462.4]
  assign _T_15490 = entriesToCheck_14_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@13464.4]
  assign _T_15491 = _T_15490 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13465.4]
  assign _T_15492 = addrQ_14 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@13466.4]
  assign conflict_14_11 = _T_15491 & _T_15492; // @[AxiLoadQueue.scala 151:68:@13467.4]
  assign _T_15494 = entriesToCheck_14_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@13469.4]
  assign _T_15495 = _T_15494 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13470.4]
  assign _T_15496 = addrQ_14 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@13471.4]
  assign conflict_14_12 = _T_15495 & _T_15496; // @[AxiLoadQueue.scala 151:68:@13472.4]
  assign _T_15498 = entriesToCheck_14_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@13474.4]
  assign _T_15499 = _T_15498 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13475.4]
  assign _T_15500 = addrQ_14 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@13476.4]
  assign conflict_14_13 = _T_15499 & _T_15500; // @[AxiLoadQueue.scala 151:68:@13477.4]
  assign _T_15502 = entriesToCheck_14_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@13479.4]
  assign _T_15503 = _T_15502 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13480.4]
  assign _T_15504 = addrQ_14 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13481.4]
  assign conflict_14_14 = _T_15503 & _T_15504; // @[AxiLoadQueue.scala 151:68:@13482.4]
  assign _T_15506 = entriesToCheck_14_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13484.4]
  assign _T_15507 = _T_15506 & addrKnown_14; // @[AxiLoadQueue.scala 151:41:@13485.4]
  assign _T_15508 = addrQ_14 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13486.4]
  assign conflict_14_15 = _T_15507 & _T_15508; // @[AxiLoadQueue.scala 151:68:@13487.4]
  assign _T_15510 = entriesToCheck_15_0 & io_storeAddrDone_0; // @[AxiLoadQueue.scala 150:92:@13489.4]
  assign _T_15511 = _T_15510 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13490.4]
  assign _T_15512 = addrQ_15 == io_storeAddrQueue_0; // @[AxiLoadQueue.scala 152:30:@13491.4]
  assign conflict_15_0 = _T_15511 & _T_15512; // @[AxiLoadQueue.scala 151:68:@13492.4]
  assign _T_15514 = entriesToCheck_15_1 & io_storeAddrDone_1; // @[AxiLoadQueue.scala 150:92:@13494.4]
  assign _T_15515 = _T_15514 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13495.4]
  assign _T_15516 = addrQ_15 == io_storeAddrQueue_1; // @[AxiLoadQueue.scala 152:30:@13496.4]
  assign conflict_15_1 = _T_15515 & _T_15516; // @[AxiLoadQueue.scala 151:68:@13497.4]
  assign _T_15518 = entriesToCheck_15_2 & io_storeAddrDone_2; // @[AxiLoadQueue.scala 150:92:@13499.4]
  assign _T_15519 = _T_15518 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13500.4]
  assign _T_15520 = addrQ_15 == io_storeAddrQueue_2; // @[AxiLoadQueue.scala 152:30:@13501.4]
  assign conflict_15_2 = _T_15519 & _T_15520; // @[AxiLoadQueue.scala 151:68:@13502.4]
  assign _T_15522 = entriesToCheck_15_3 & io_storeAddrDone_3; // @[AxiLoadQueue.scala 150:92:@13504.4]
  assign _T_15523 = _T_15522 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13505.4]
  assign _T_15524 = addrQ_15 == io_storeAddrQueue_3; // @[AxiLoadQueue.scala 152:30:@13506.4]
  assign conflict_15_3 = _T_15523 & _T_15524; // @[AxiLoadQueue.scala 151:68:@13507.4]
  assign _T_15526 = entriesToCheck_15_4 & io_storeAddrDone_4; // @[AxiLoadQueue.scala 150:92:@13509.4]
  assign _T_15527 = _T_15526 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13510.4]
  assign _T_15528 = addrQ_15 == io_storeAddrQueue_4; // @[AxiLoadQueue.scala 152:30:@13511.4]
  assign conflict_15_4 = _T_15527 & _T_15528; // @[AxiLoadQueue.scala 151:68:@13512.4]
  assign _T_15530 = entriesToCheck_15_5 & io_storeAddrDone_5; // @[AxiLoadQueue.scala 150:92:@13514.4]
  assign _T_15531 = _T_15530 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13515.4]
  assign _T_15532 = addrQ_15 == io_storeAddrQueue_5; // @[AxiLoadQueue.scala 152:30:@13516.4]
  assign conflict_15_5 = _T_15531 & _T_15532; // @[AxiLoadQueue.scala 151:68:@13517.4]
  assign _T_15534 = entriesToCheck_15_6 & io_storeAddrDone_6; // @[AxiLoadQueue.scala 150:92:@13519.4]
  assign _T_15535 = _T_15534 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13520.4]
  assign _T_15536 = addrQ_15 == io_storeAddrQueue_6; // @[AxiLoadQueue.scala 152:30:@13521.4]
  assign conflict_15_6 = _T_15535 & _T_15536; // @[AxiLoadQueue.scala 151:68:@13522.4]
  assign _T_15538 = entriesToCheck_15_7 & io_storeAddrDone_7; // @[AxiLoadQueue.scala 150:92:@13524.4]
  assign _T_15539 = _T_15538 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13525.4]
  assign _T_15540 = addrQ_15 == io_storeAddrQueue_7; // @[AxiLoadQueue.scala 152:30:@13526.4]
  assign conflict_15_7 = _T_15539 & _T_15540; // @[AxiLoadQueue.scala 151:68:@13527.4]
  assign _T_15542 = entriesToCheck_15_8 & io_storeAddrDone_8; // @[AxiLoadQueue.scala 150:92:@13529.4]
  assign _T_15543 = _T_15542 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13530.4]
  assign _T_15544 = addrQ_15 == io_storeAddrQueue_8; // @[AxiLoadQueue.scala 152:30:@13531.4]
  assign conflict_15_8 = _T_15543 & _T_15544; // @[AxiLoadQueue.scala 151:68:@13532.4]
  assign _T_15546 = entriesToCheck_15_9 & io_storeAddrDone_9; // @[AxiLoadQueue.scala 150:92:@13534.4]
  assign _T_15547 = _T_15546 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13535.4]
  assign _T_15548 = addrQ_15 == io_storeAddrQueue_9; // @[AxiLoadQueue.scala 152:30:@13536.4]
  assign conflict_15_9 = _T_15547 & _T_15548; // @[AxiLoadQueue.scala 151:68:@13537.4]
  assign _T_15550 = entriesToCheck_15_10 & io_storeAddrDone_10; // @[AxiLoadQueue.scala 150:92:@13539.4]
  assign _T_15551 = _T_15550 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13540.4]
  assign _T_15552 = addrQ_15 == io_storeAddrQueue_10; // @[AxiLoadQueue.scala 152:30:@13541.4]
  assign conflict_15_10 = _T_15551 & _T_15552; // @[AxiLoadQueue.scala 151:68:@13542.4]
  assign _T_15554 = entriesToCheck_15_11 & io_storeAddrDone_11; // @[AxiLoadQueue.scala 150:92:@13544.4]
  assign _T_15555 = _T_15554 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13545.4]
  assign _T_15556 = addrQ_15 == io_storeAddrQueue_11; // @[AxiLoadQueue.scala 152:30:@13546.4]
  assign conflict_15_11 = _T_15555 & _T_15556; // @[AxiLoadQueue.scala 151:68:@13547.4]
  assign _T_15558 = entriesToCheck_15_12 & io_storeAddrDone_12; // @[AxiLoadQueue.scala 150:92:@13549.4]
  assign _T_15559 = _T_15558 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13550.4]
  assign _T_15560 = addrQ_15 == io_storeAddrQueue_12; // @[AxiLoadQueue.scala 152:30:@13551.4]
  assign conflict_15_12 = _T_15559 & _T_15560; // @[AxiLoadQueue.scala 151:68:@13552.4]
  assign _T_15562 = entriesToCheck_15_13 & io_storeAddrDone_13; // @[AxiLoadQueue.scala 150:92:@13554.4]
  assign _T_15563 = _T_15562 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13555.4]
  assign _T_15564 = addrQ_15 == io_storeAddrQueue_13; // @[AxiLoadQueue.scala 152:30:@13556.4]
  assign conflict_15_13 = _T_15563 & _T_15564; // @[AxiLoadQueue.scala 151:68:@13557.4]
  assign _T_15566 = entriesToCheck_15_14 & io_storeAddrDone_14; // @[AxiLoadQueue.scala 150:92:@13559.4]
  assign _T_15567 = _T_15566 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13560.4]
  assign _T_15568 = addrQ_15 == io_storeAddrQueue_14; // @[AxiLoadQueue.scala 152:30:@13561.4]
  assign conflict_15_14 = _T_15567 & _T_15568; // @[AxiLoadQueue.scala 151:68:@13562.4]
  assign _T_15570 = entriesToCheck_15_15 & io_storeAddrDone_15; // @[AxiLoadQueue.scala 150:92:@13564.4]
  assign _T_15571 = _T_15570 & addrKnown_15; // @[AxiLoadQueue.scala 151:41:@13565.4]
  assign _T_15572 = addrQ_15 == io_storeAddrQueue_15; // @[AxiLoadQueue.scala 152:30:@13566.4]
  assign conflict_15_15 = _T_15571 & _T_15572; // @[AxiLoadQueue.scala 151:68:@13567.4]
  assign _T_16805 = io_storeAddrDone_0 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13570.4]
  assign storeAddrNotKnownFlags_0_0 = _T_16805 & entriesToCheck_0_0; // @[AxiLoadQueue.scala 163:19:@13571.4]
  assign _T_16808 = io_storeAddrDone_1 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13572.4]
  assign storeAddrNotKnownFlags_0_1 = _T_16808 & entriesToCheck_0_1; // @[AxiLoadQueue.scala 163:19:@13573.4]
  assign _T_16811 = io_storeAddrDone_2 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13574.4]
  assign storeAddrNotKnownFlags_0_2 = _T_16811 & entriesToCheck_0_2; // @[AxiLoadQueue.scala 163:19:@13575.4]
  assign _T_16814 = io_storeAddrDone_3 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13576.4]
  assign storeAddrNotKnownFlags_0_3 = _T_16814 & entriesToCheck_0_3; // @[AxiLoadQueue.scala 163:19:@13577.4]
  assign _T_16817 = io_storeAddrDone_4 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13578.4]
  assign storeAddrNotKnownFlags_0_4 = _T_16817 & entriesToCheck_0_4; // @[AxiLoadQueue.scala 163:19:@13579.4]
  assign _T_16820 = io_storeAddrDone_5 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13580.4]
  assign storeAddrNotKnownFlags_0_5 = _T_16820 & entriesToCheck_0_5; // @[AxiLoadQueue.scala 163:19:@13581.4]
  assign _T_16823 = io_storeAddrDone_6 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13582.4]
  assign storeAddrNotKnownFlags_0_6 = _T_16823 & entriesToCheck_0_6; // @[AxiLoadQueue.scala 163:19:@13583.4]
  assign _T_16826 = io_storeAddrDone_7 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13584.4]
  assign storeAddrNotKnownFlags_0_7 = _T_16826 & entriesToCheck_0_7; // @[AxiLoadQueue.scala 163:19:@13585.4]
  assign _T_16829 = io_storeAddrDone_8 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13586.4]
  assign storeAddrNotKnownFlags_0_8 = _T_16829 & entriesToCheck_0_8; // @[AxiLoadQueue.scala 163:19:@13587.4]
  assign _T_16832 = io_storeAddrDone_9 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13588.4]
  assign storeAddrNotKnownFlags_0_9 = _T_16832 & entriesToCheck_0_9; // @[AxiLoadQueue.scala 163:19:@13589.4]
  assign _T_16835 = io_storeAddrDone_10 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13590.4]
  assign storeAddrNotKnownFlags_0_10 = _T_16835 & entriesToCheck_0_10; // @[AxiLoadQueue.scala 163:19:@13591.4]
  assign _T_16838 = io_storeAddrDone_11 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13592.4]
  assign storeAddrNotKnownFlags_0_11 = _T_16838 & entriesToCheck_0_11; // @[AxiLoadQueue.scala 163:19:@13593.4]
  assign _T_16841 = io_storeAddrDone_12 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13594.4]
  assign storeAddrNotKnownFlags_0_12 = _T_16841 & entriesToCheck_0_12; // @[AxiLoadQueue.scala 163:19:@13595.4]
  assign _T_16844 = io_storeAddrDone_13 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13596.4]
  assign storeAddrNotKnownFlags_0_13 = _T_16844 & entriesToCheck_0_13; // @[AxiLoadQueue.scala 163:19:@13597.4]
  assign _T_16847 = io_storeAddrDone_14 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13598.4]
  assign storeAddrNotKnownFlags_0_14 = _T_16847 & entriesToCheck_0_14; // @[AxiLoadQueue.scala 163:19:@13599.4]
  assign _T_16850 = io_storeAddrDone_15 == 1'h0; // @[AxiLoadQueue.scala 163:13:@13600.4]
  assign storeAddrNotKnownFlags_0_15 = _T_16850 & entriesToCheck_0_15; // @[AxiLoadQueue.scala 163:19:@13601.4]
  assign storeAddrNotKnownFlags_1_0 = _T_16805 & entriesToCheck_1_0; // @[AxiLoadQueue.scala 163:19:@13619.4]
  assign storeAddrNotKnownFlags_1_1 = _T_16808 & entriesToCheck_1_1; // @[AxiLoadQueue.scala 163:19:@13621.4]
  assign storeAddrNotKnownFlags_1_2 = _T_16811 & entriesToCheck_1_2; // @[AxiLoadQueue.scala 163:19:@13623.4]
  assign storeAddrNotKnownFlags_1_3 = _T_16814 & entriesToCheck_1_3; // @[AxiLoadQueue.scala 163:19:@13625.4]
  assign storeAddrNotKnownFlags_1_4 = _T_16817 & entriesToCheck_1_4; // @[AxiLoadQueue.scala 163:19:@13627.4]
  assign storeAddrNotKnownFlags_1_5 = _T_16820 & entriesToCheck_1_5; // @[AxiLoadQueue.scala 163:19:@13629.4]
  assign storeAddrNotKnownFlags_1_6 = _T_16823 & entriesToCheck_1_6; // @[AxiLoadQueue.scala 163:19:@13631.4]
  assign storeAddrNotKnownFlags_1_7 = _T_16826 & entriesToCheck_1_7; // @[AxiLoadQueue.scala 163:19:@13633.4]
  assign storeAddrNotKnownFlags_1_8 = _T_16829 & entriesToCheck_1_8; // @[AxiLoadQueue.scala 163:19:@13635.4]
  assign storeAddrNotKnownFlags_1_9 = _T_16832 & entriesToCheck_1_9; // @[AxiLoadQueue.scala 163:19:@13637.4]
  assign storeAddrNotKnownFlags_1_10 = _T_16835 & entriesToCheck_1_10; // @[AxiLoadQueue.scala 163:19:@13639.4]
  assign storeAddrNotKnownFlags_1_11 = _T_16838 & entriesToCheck_1_11; // @[AxiLoadQueue.scala 163:19:@13641.4]
  assign storeAddrNotKnownFlags_1_12 = _T_16841 & entriesToCheck_1_12; // @[AxiLoadQueue.scala 163:19:@13643.4]
  assign storeAddrNotKnownFlags_1_13 = _T_16844 & entriesToCheck_1_13; // @[AxiLoadQueue.scala 163:19:@13645.4]
  assign storeAddrNotKnownFlags_1_14 = _T_16847 & entriesToCheck_1_14; // @[AxiLoadQueue.scala 163:19:@13647.4]
  assign storeAddrNotKnownFlags_1_15 = _T_16850 & entriesToCheck_1_15; // @[AxiLoadQueue.scala 163:19:@13649.4]
  assign storeAddrNotKnownFlags_2_0 = _T_16805 & entriesToCheck_2_0; // @[AxiLoadQueue.scala 163:19:@13667.4]
  assign storeAddrNotKnownFlags_2_1 = _T_16808 & entriesToCheck_2_1; // @[AxiLoadQueue.scala 163:19:@13669.4]
  assign storeAddrNotKnownFlags_2_2 = _T_16811 & entriesToCheck_2_2; // @[AxiLoadQueue.scala 163:19:@13671.4]
  assign storeAddrNotKnownFlags_2_3 = _T_16814 & entriesToCheck_2_3; // @[AxiLoadQueue.scala 163:19:@13673.4]
  assign storeAddrNotKnownFlags_2_4 = _T_16817 & entriesToCheck_2_4; // @[AxiLoadQueue.scala 163:19:@13675.4]
  assign storeAddrNotKnownFlags_2_5 = _T_16820 & entriesToCheck_2_5; // @[AxiLoadQueue.scala 163:19:@13677.4]
  assign storeAddrNotKnownFlags_2_6 = _T_16823 & entriesToCheck_2_6; // @[AxiLoadQueue.scala 163:19:@13679.4]
  assign storeAddrNotKnownFlags_2_7 = _T_16826 & entriesToCheck_2_7; // @[AxiLoadQueue.scala 163:19:@13681.4]
  assign storeAddrNotKnownFlags_2_8 = _T_16829 & entriesToCheck_2_8; // @[AxiLoadQueue.scala 163:19:@13683.4]
  assign storeAddrNotKnownFlags_2_9 = _T_16832 & entriesToCheck_2_9; // @[AxiLoadQueue.scala 163:19:@13685.4]
  assign storeAddrNotKnownFlags_2_10 = _T_16835 & entriesToCheck_2_10; // @[AxiLoadQueue.scala 163:19:@13687.4]
  assign storeAddrNotKnownFlags_2_11 = _T_16838 & entriesToCheck_2_11; // @[AxiLoadQueue.scala 163:19:@13689.4]
  assign storeAddrNotKnownFlags_2_12 = _T_16841 & entriesToCheck_2_12; // @[AxiLoadQueue.scala 163:19:@13691.4]
  assign storeAddrNotKnownFlags_2_13 = _T_16844 & entriesToCheck_2_13; // @[AxiLoadQueue.scala 163:19:@13693.4]
  assign storeAddrNotKnownFlags_2_14 = _T_16847 & entriesToCheck_2_14; // @[AxiLoadQueue.scala 163:19:@13695.4]
  assign storeAddrNotKnownFlags_2_15 = _T_16850 & entriesToCheck_2_15; // @[AxiLoadQueue.scala 163:19:@13697.4]
  assign storeAddrNotKnownFlags_3_0 = _T_16805 & entriesToCheck_3_0; // @[AxiLoadQueue.scala 163:19:@13715.4]
  assign storeAddrNotKnownFlags_3_1 = _T_16808 & entriesToCheck_3_1; // @[AxiLoadQueue.scala 163:19:@13717.4]
  assign storeAddrNotKnownFlags_3_2 = _T_16811 & entriesToCheck_3_2; // @[AxiLoadQueue.scala 163:19:@13719.4]
  assign storeAddrNotKnownFlags_3_3 = _T_16814 & entriesToCheck_3_3; // @[AxiLoadQueue.scala 163:19:@13721.4]
  assign storeAddrNotKnownFlags_3_4 = _T_16817 & entriesToCheck_3_4; // @[AxiLoadQueue.scala 163:19:@13723.4]
  assign storeAddrNotKnownFlags_3_5 = _T_16820 & entriesToCheck_3_5; // @[AxiLoadQueue.scala 163:19:@13725.4]
  assign storeAddrNotKnownFlags_3_6 = _T_16823 & entriesToCheck_3_6; // @[AxiLoadQueue.scala 163:19:@13727.4]
  assign storeAddrNotKnownFlags_3_7 = _T_16826 & entriesToCheck_3_7; // @[AxiLoadQueue.scala 163:19:@13729.4]
  assign storeAddrNotKnownFlags_3_8 = _T_16829 & entriesToCheck_3_8; // @[AxiLoadQueue.scala 163:19:@13731.4]
  assign storeAddrNotKnownFlags_3_9 = _T_16832 & entriesToCheck_3_9; // @[AxiLoadQueue.scala 163:19:@13733.4]
  assign storeAddrNotKnownFlags_3_10 = _T_16835 & entriesToCheck_3_10; // @[AxiLoadQueue.scala 163:19:@13735.4]
  assign storeAddrNotKnownFlags_3_11 = _T_16838 & entriesToCheck_3_11; // @[AxiLoadQueue.scala 163:19:@13737.4]
  assign storeAddrNotKnownFlags_3_12 = _T_16841 & entriesToCheck_3_12; // @[AxiLoadQueue.scala 163:19:@13739.4]
  assign storeAddrNotKnownFlags_3_13 = _T_16844 & entriesToCheck_3_13; // @[AxiLoadQueue.scala 163:19:@13741.4]
  assign storeAddrNotKnownFlags_3_14 = _T_16847 & entriesToCheck_3_14; // @[AxiLoadQueue.scala 163:19:@13743.4]
  assign storeAddrNotKnownFlags_3_15 = _T_16850 & entriesToCheck_3_15; // @[AxiLoadQueue.scala 163:19:@13745.4]
  assign storeAddrNotKnownFlags_4_0 = _T_16805 & entriesToCheck_4_0; // @[AxiLoadQueue.scala 163:19:@13763.4]
  assign storeAddrNotKnownFlags_4_1 = _T_16808 & entriesToCheck_4_1; // @[AxiLoadQueue.scala 163:19:@13765.4]
  assign storeAddrNotKnownFlags_4_2 = _T_16811 & entriesToCheck_4_2; // @[AxiLoadQueue.scala 163:19:@13767.4]
  assign storeAddrNotKnownFlags_4_3 = _T_16814 & entriesToCheck_4_3; // @[AxiLoadQueue.scala 163:19:@13769.4]
  assign storeAddrNotKnownFlags_4_4 = _T_16817 & entriesToCheck_4_4; // @[AxiLoadQueue.scala 163:19:@13771.4]
  assign storeAddrNotKnownFlags_4_5 = _T_16820 & entriesToCheck_4_5; // @[AxiLoadQueue.scala 163:19:@13773.4]
  assign storeAddrNotKnownFlags_4_6 = _T_16823 & entriesToCheck_4_6; // @[AxiLoadQueue.scala 163:19:@13775.4]
  assign storeAddrNotKnownFlags_4_7 = _T_16826 & entriesToCheck_4_7; // @[AxiLoadQueue.scala 163:19:@13777.4]
  assign storeAddrNotKnownFlags_4_8 = _T_16829 & entriesToCheck_4_8; // @[AxiLoadQueue.scala 163:19:@13779.4]
  assign storeAddrNotKnownFlags_4_9 = _T_16832 & entriesToCheck_4_9; // @[AxiLoadQueue.scala 163:19:@13781.4]
  assign storeAddrNotKnownFlags_4_10 = _T_16835 & entriesToCheck_4_10; // @[AxiLoadQueue.scala 163:19:@13783.4]
  assign storeAddrNotKnownFlags_4_11 = _T_16838 & entriesToCheck_4_11; // @[AxiLoadQueue.scala 163:19:@13785.4]
  assign storeAddrNotKnownFlags_4_12 = _T_16841 & entriesToCheck_4_12; // @[AxiLoadQueue.scala 163:19:@13787.4]
  assign storeAddrNotKnownFlags_4_13 = _T_16844 & entriesToCheck_4_13; // @[AxiLoadQueue.scala 163:19:@13789.4]
  assign storeAddrNotKnownFlags_4_14 = _T_16847 & entriesToCheck_4_14; // @[AxiLoadQueue.scala 163:19:@13791.4]
  assign storeAddrNotKnownFlags_4_15 = _T_16850 & entriesToCheck_4_15; // @[AxiLoadQueue.scala 163:19:@13793.4]
  assign storeAddrNotKnownFlags_5_0 = _T_16805 & entriesToCheck_5_0; // @[AxiLoadQueue.scala 163:19:@13811.4]
  assign storeAddrNotKnownFlags_5_1 = _T_16808 & entriesToCheck_5_1; // @[AxiLoadQueue.scala 163:19:@13813.4]
  assign storeAddrNotKnownFlags_5_2 = _T_16811 & entriesToCheck_5_2; // @[AxiLoadQueue.scala 163:19:@13815.4]
  assign storeAddrNotKnownFlags_5_3 = _T_16814 & entriesToCheck_5_3; // @[AxiLoadQueue.scala 163:19:@13817.4]
  assign storeAddrNotKnownFlags_5_4 = _T_16817 & entriesToCheck_5_4; // @[AxiLoadQueue.scala 163:19:@13819.4]
  assign storeAddrNotKnownFlags_5_5 = _T_16820 & entriesToCheck_5_5; // @[AxiLoadQueue.scala 163:19:@13821.4]
  assign storeAddrNotKnownFlags_5_6 = _T_16823 & entriesToCheck_5_6; // @[AxiLoadQueue.scala 163:19:@13823.4]
  assign storeAddrNotKnownFlags_5_7 = _T_16826 & entriesToCheck_5_7; // @[AxiLoadQueue.scala 163:19:@13825.4]
  assign storeAddrNotKnownFlags_5_8 = _T_16829 & entriesToCheck_5_8; // @[AxiLoadQueue.scala 163:19:@13827.4]
  assign storeAddrNotKnownFlags_5_9 = _T_16832 & entriesToCheck_5_9; // @[AxiLoadQueue.scala 163:19:@13829.4]
  assign storeAddrNotKnownFlags_5_10 = _T_16835 & entriesToCheck_5_10; // @[AxiLoadQueue.scala 163:19:@13831.4]
  assign storeAddrNotKnownFlags_5_11 = _T_16838 & entriesToCheck_5_11; // @[AxiLoadQueue.scala 163:19:@13833.4]
  assign storeAddrNotKnownFlags_5_12 = _T_16841 & entriesToCheck_5_12; // @[AxiLoadQueue.scala 163:19:@13835.4]
  assign storeAddrNotKnownFlags_5_13 = _T_16844 & entriesToCheck_5_13; // @[AxiLoadQueue.scala 163:19:@13837.4]
  assign storeAddrNotKnownFlags_5_14 = _T_16847 & entriesToCheck_5_14; // @[AxiLoadQueue.scala 163:19:@13839.4]
  assign storeAddrNotKnownFlags_5_15 = _T_16850 & entriesToCheck_5_15; // @[AxiLoadQueue.scala 163:19:@13841.4]
  assign storeAddrNotKnownFlags_6_0 = _T_16805 & entriesToCheck_6_0; // @[AxiLoadQueue.scala 163:19:@13859.4]
  assign storeAddrNotKnownFlags_6_1 = _T_16808 & entriesToCheck_6_1; // @[AxiLoadQueue.scala 163:19:@13861.4]
  assign storeAddrNotKnownFlags_6_2 = _T_16811 & entriesToCheck_6_2; // @[AxiLoadQueue.scala 163:19:@13863.4]
  assign storeAddrNotKnownFlags_6_3 = _T_16814 & entriesToCheck_6_3; // @[AxiLoadQueue.scala 163:19:@13865.4]
  assign storeAddrNotKnownFlags_6_4 = _T_16817 & entriesToCheck_6_4; // @[AxiLoadQueue.scala 163:19:@13867.4]
  assign storeAddrNotKnownFlags_6_5 = _T_16820 & entriesToCheck_6_5; // @[AxiLoadQueue.scala 163:19:@13869.4]
  assign storeAddrNotKnownFlags_6_6 = _T_16823 & entriesToCheck_6_6; // @[AxiLoadQueue.scala 163:19:@13871.4]
  assign storeAddrNotKnownFlags_6_7 = _T_16826 & entriesToCheck_6_7; // @[AxiLoadQueue.scala 163:19:@13873.4]
  assign storeAddrNotKnownFlags_6_8 = _T_16829 & entriesToCheck_6_8; // @[AxiLoadQueue.scala 163:19:@13875.4]
  assign storeAddrNotKnownFlags_6_9 = _T_16832 & entriesToCheck_6_9; // @[AxiLoadQueue.scala 163:19:@13877.4]
  assign storeAddrNotKnownFlags_6_10 = _T_16835 & entriesToCheck_6_10; // @[AxiLoadQueue.scala 163:19:@13879.4]
  assign storeAddrNotKnownFlags_6_11 = _T_16838 & entriesToCheck_6_11; // @[AxiLoadQueue.scala 163:19:@13881.4]
  assign storeAddrNotKnownFlags_6_12 = _T_16841 & entriesToCheck_6_12; // @[AxiLoadQueue.scala 163:19:@13883.4]
  assign storeAddrNotKnownFlags_6_13 = _T_16844 & entriesToCheck_6_13; // @[AxiLoadQueue.scala 163:19:@13885.4]
  assign storeAddrNotKnownFlags_6_14 = _T_16847 & entriesToCheck_6_14; // @[AxiLoadQueue.scala 163:19:@13887.4]
  assign storeAddrNotKnownFlags_6_15 = _T_16850 & entriesToCheck_6_15; // @[AxiLoadQueue.scala 163:19:@13889.4]
  assign storeAddrNotKnownFlags_7_0 = _T_16805 & entriesToCheck_7_0; // @[AxiLoadQueue.scala 163:19:@13907.4]
  assign storeAddrNotKnownFlags_7_1 = _T_16808 & entriesToCheck_7_1; // @[AxiLoadQueue.scala 163:19:@13909.4]
  assign storeAddrNotKnownFlags_7_2 = _T_16811 & entriesToCheck_7_2; // @[AxiLoadQueue.scala 163:19:@13911.4]
  assign storeAddrNotKnownFlags_7_3 = _T_16814 & entriesToCheck_7_3; // @[AxiLoadQueue.scala 163:19:@13913.4]
  assign storeAddrNotKnownFlags_7_4 = _T_16817 & entriesToCheck_7_4; // @[AxiLoadQueue.scala 163:19:@13915.4]
  assign storeAddrNotKnownFlags_7_5 = _T_16820 & entriesToCheck_7_5; // @[AxiLoadQueue.scala 163:19:@13917.4]
  assign storeAddrNotKnownFlags_7_6 = _T_16823 & entriesToCheck_7_6; // @[AxiLoadQueue.scala 163:19:@13919.4]
  assign storeAddrNotKnownFlags_7_7 = _T_16826 & entriesToCheck_7_7; // @[AxiLoadQueue.scala 163:19:@13921.4]
  assign storeAddrNotKnownFlags_7_8 = _T_16829 & entriesToCheck_7_8; // @[AxiLoadQueue.scala 163:19:@13923.4]
  assign storeAddrNotKnownFlags_7_9 = _T_16832 & entriesToCheck_7_9; // @[AxiLoadQueue.scala 163:19:@13925.4]
  assign storeAddrNotKnownFlags_7_10 = _T_16835 & entriesToCheck_7_10; // @[AxiLoadQueue.scala 163:19:@13927.4]
  assign storeAddrNotKnownFlags_7_11 = _T_16838 & entriesToCheck_7_11; // @[AxiLoadQueue.scala 163:19:@13929.4]
  assign storeAddrNotKnownFlags_7_12 = _T_16841 & entriesToCheck_7_12; // @[AxiLoadQueue.scala 163:19:@13931.4]
  assign storeAddrNotKnownFlags_7_13 = _T_16844 & entriesToCheck_7_13; // @[AxiLoadQueue.scala 163:19:@13933.4]
  assign storeAddrNotKnownFlags_7_14 = _T_16847 & entriesToCheck_7_14; // @[AxiLoadQueue.scala 163:19:@13935.4]
  assign storeAddrNotKnownFlags_7_15 = _T_16850 & entriesToCheck_7_15; // @[AxiLoadQueue.scala 163:19:@13937.4]
  assign storeAddrNotKnownFlags_8_0 = _T_16805 & entriesToCheck_8_0; // @[AxiLoadQueue.scala 163:19:@13955.4]
  assign storeAddrNotKnownFlags_8_1 = _T_16808 & entriesToCheck_8_1; // @[AxiLoadQueue.scala 163:19:@13957.4]
  assign storeAddrNotKnownFlags_8_2 = _T_16811 & entriesToCheck_8_2; // @[AxiLoadQueue.scala 163:19:@13959.4]
  assign storeAddrNotKnownFlags_8_3 = _T_16814 & entriesToCheck_8_3; // @[AxiLoadQueue.scala 163:19:@13961.4]
  assign storeAddrNotKnownFlags_8_4 = _T_16817 & entriesToCheck_8_4; // @[AxiLoadQueue.scala 163:19:@13963.4]
  assign storeAddrNotKnownFlags_8_5 = _T_16820 & entriesToCheck_8_5; // @[AxiLoadQueue.scala 163:19:@13965.4]
  assign storeAddrNotKnownFlags_8_6 = _T_16823 & entriesToCheck_8_6; // @[AxiLoadQueue.scala 163:19:@13967.4]
  assign storeAddrNotKnownFlags_8_7 = _T_16826 & entriesToCheck_8_7; // @[AxiLoadQueue.scala 163:19:@13969.4]
  assign storeAddrNotKnownFlags_8_8 = _T_16829 & entriesToCheck_8_8; // @[AxiLoadQueue.scala 163:19:@13971.4]
  assign storeAddrNotKnownFlags_8_9 = _T_16832 & entriesToCheck_8_9; // @[AxiLoadQueue.scala 163:19:@13973.4]
  assign storeAddrNotKnownFlags_8_10 = _T_16835 & entriesToCheck_8_10; // @[AxiLoadQueue.scala 163:19:@13975.4]
  assign storeAddrNotKnownFlags_8_11 = _T_16838 & entriesToCheck_8_11; // @[AxiLoadQueue.scala 163:19:@13977.4]
  assign storeAddrNotKnownFlags_8_12 = _T_16841 & entriesToCheck_8_12; // @[AxiLoadQueue.scala 163:19:@13979.4]
  assign storeAddrNotKnownFlags_8_13 = _T_16844 & entriesToCheck_8_13; // @[AxiLoadQueue.scala 163:19:@13981.4]
  assign storeAddrNotKnownFlags_8_14 = _T_16847 & entriesToCheck_8_14; // @[AxiLoadQueue.scala 163:19:@13983.4]
  assign storeAddrNotKnownFlags_8_15 = _T_16850 & entriesToCheck_8_15; // @[AxiLoadQueue.scala 163:19:@13985.4]
  assign storeAddrNotKnownFlags_9_0 = _T_16805 & entriesToCheck_9_0; // @[AxiLoadQueue.scala 163:19:@14003.4]
  assign storeAddrNotKnownFlags_9_1 = _T_16808 & entriesToCheck_9_1; // @[AxiLoadQueue.scala 163:19:@14005.4]
  assign storeAddrNotKnownFlags_9_2 = _T_16811 & entriesToCheck_9_2; // @[AxiLoadQueue.scala 163:19:@14007.4]
  assign storeAddrNotKnownFlags_9_3 = _T_16814 & entriesToCheck_9_3; // @[AxiLoadQueue.scala 163:19:@14009.4]
  assign storeAddrNotKnownFlags_9_4 = _T_16817 & entriesToCheck_9_4; // @[AxiLoadQueue.scala 163:19:@14011.4]
  assign storeAddrNotKnownFlags_9_5 = _T_16820 & entriesToCheck_9_5; // @[AxiLoadQueue.scala 163:19:@14013.4]
  assign storeAddrNotKnownFlags_9_6 = _T_16823 & entriesToCheck_9_6; // @[AxiLoadQueue.scala 163:19:@14015.4]
  assign storeAddrNotKnownFlags_9_7 = _T_16826 & entriesToCheck_9_7; // @[AxiLoadQueue.scala 163:19:@14017.4]
  assign storeAddrNotKnownFlags_9_8 = _T_16829 & entriesToCheck_9_8; // @[AxiLoadQueue.scala 163:19:@14019.4]
  assign storeAddrNotKnownFlags_9_9 = _T_16832 & entriesToCheck_9_9; // @[AxiLoadQueue.scala 163:19:@14021.4]
  assign storeAddrNotKnownFlags_9_10 = _T_16835 & entriesToCheck_9_10; // @[AxiLoadQueue.scala 163:19:@14023.4]
  assign storeAddrNotKnownFlags_9_11 = _T_16838 & entriesToCheck_9_11; // @[AxiLoadQueue.scala 163:19:@14025.4]
  assign storeAddrNotKnownFlags_9_12 = _T_16841 & entriesToCheck_9_12; // @[AxiLoadQueue.scala 163:19:@14027.4]
  assign storeAddrNotKnownFlags_9_13 = _T_16844 & entriesToCheck_9_13; // @[AxiLoadQueue.scala 163:19:@14029.4]
  assign storeAddrNotKnownFlags_9_14 = _T_16847 & entriesToCheck_9_14; // @[AxiLoadQueue.scala 163:19:@14031.4]
  assign storeAddrNotKnownFlags_9_15 = _T_16850 & entriesToCheck_9_15; // @[AxiLoadQueue.scala 163:19:@14033.4]
  assign storeAddrNotKnownFlags_10_0 = _T_16805 & entriesToCheck_10_0; // @[AxiLoadQueue.scala 163:19:@14051.4]
  assign storeAddrNotKnownFlags_10_1 = _T_16808 & entriesToCheck_10_1; // @[AxiLoadQueue.scala 163:19:@14053.4]
  assign storeAddrNotKnownFlags_10_2 = _T_16811 & entriesToCheck_10_2; // @[AxiLoadQueue.scala 163:19:@14055.4]
  assign storeAddrNotKnownFlags_10_3 = _T_16814 & entriesToCheck_10_3; // @[AxiLoadQueue.scala 163:19:@14057.4]
  assign storeAddrNotKnownFlags_10_4 = _T_16817 & entriesToCheck_10_4; // @[AxiLoadQueue.scala 163:19:@14059.4]
  assign storeAddrNotKnownFlags_10_5 = _T_16820 & entriesToCheck_10_5; // @[AxiLoadQueue.scala 163:19:@14061.4]
  assign storeAddrNotKnownFlags_10_6 = _T_16823 & entriesToCheck_10_6; // @[AxiLoadQueue.scala 163:19:@14063.4]
  assign storeAddrNotKnownFlags_10_7 = _T_16826 & entriesToCheck_10_7; // @[AxiLoadQueue.scala 163:19:@14065.4]
  assign storeAddrNotKnownFlags_10_8 = _T_16829 & entriesToCheck_10_8; // @[AxiLoadQueue.scala 163:19:@14067.4]
  assign storeAddrNotKnownFlags_10_9 = _T_16832 & entriesToCheck_10_9; // @[AxiLoadQueue.scala 163:19:@14069.4]
  assign storeAddrNotKnownFlags_10_10 = _T_16835 & entriesToCheck_10_10; // @[AxiLoadQueue.scala 163:19:@14071.4]
  assign storeAddrNotKnownFlags_10_11 = _T_16838 & entriesToCheck_10_11; // @[AxiLoadQueue.scala 163:19:@14073.4]
  assign storeAddrNotKnownFlags_10_12 = _T_16841 & entriesToCheck_10_12; // @[AxiLoadQueue.scala 163:19:@14075.4]
  assign storeAddrNotKnownFlags_10_13 = _T_16844 & entriesToCheck_10_13; // @[AxiLoadQueue.scala 163:19:@14077.4]
  assign storeAddrNotKnownFlags_10_14 = _T_16847 & entriesToCheck_10_14; // @[AxiLoadQueue.scala 163:19:@14079.4]
  assign storeAddrNotKnownFlags_10_15 = _T_16850 & entriesToCheck_10_15; // @[AxiLoadQueue.scala 163:19:@14081.4]
  assign storeAddrNotKnownFlags_11_0 = _T_16805 & entriesToCheck_11_0; // @[AxiLoadQueue.scala 163:19:@14099.4]
  assign storeAddrNotKnownFlags_11_1 = _T_16808 & entriesToCheck_11_1; // @[AxiLoadQueue.scala 163:19:@14101.4]
  assign storeAddrNotKnownFlags_11_2 = _T_16811 & entriesToCheck_11_2; // @[AxiLoadQueue.scala 163:19:@14103.4]
  assign storeAddrNotKnownFlags_11_3 = _T_16814 & entriesToCheck_11_3; // @[AxiLoadQueue.scala 163:19:@14105.4]
  assign storeAddrNotKnownFlags_11_4 = _T_16817 & entriesToCheck_11_4; // @[AxiLoadQueue.scala 163:19:@14107.4]
  assign storeAddrNotKnownFlags_11_5 = _T_16820 & entriesToCheck_11_5; // @[AxiLoadQueue.scala 163:19:@14109.4]
  assign storeAddrNotKnownFlags_11_6 = _T_16823 & entriesToCheck_11_6; // @[AxiLoadQueue.scala 163:19:@14111.4]
  assign storeAddrNotKnownFlags_11_7 = _T_16826 & entriesToCheck_11_7; // @[AxiLoadQueue.scala 163:19:@14113.4]
  assign storeAddrNotKnownFlags_11_8 = _T_16829 & entriesToCheck_11_8; // @[AxiLoadQueue.scala 163:19:@14115.4]
  assign storeAddrNotKnownFlags_11_9 = _T_16832 & entriesToCheck_11_9; // @[AxiLoadQueue.scala 163:19:@14117.4]
  assign storeAddrNotKnownFlags_11_10 = _T_16835 & entriesToCheck_11_10; // @[AxiLoadQueue.scala 163:19:@14119.4]
  assign storeAddrNotKnownFlags_11_11 = _T_16838 & entriesToCheck_11_11; // @[AxiLoadQueue.scala 163:19:@14121.4]
  assign storeAddrNotKnownFlags_11_12 = _T_16841 & entriesToCheck_11_12; // @[AxiLoadQueue.scala 163:19:@14123.4]
  assign storeAddrNotKnownFlags_11_13 = _T_16844 & entriesToCheck_11_13; // @[AxiLoadQueue.scala 163:19:@14125.4]
  assign storeAddrNotKnownFlags_11_14 = _T_16847 & entriesToCheck_11_14; // @[AxiLoadQueue.scala 163:19:@14127.4]
  assign storeAddrNotKnownFlags_11_15 = _T_16850 & entriesToCheck_11_15; // @[AxiLoadQueue.scala 163:19:@14129.4]
  assign storeAddrNotKnownFlags_12_0 = _T_16805 & entriesToCheck_12_0; // @[AxiLoadQueue.scala 163:19:@14147.4]
  assign storeAddrNotKnownFlags_12_1 = _T_16808 & entriesToCheck_12_1; // @[AxiLoadQueue.scala 163:19:@14149.4]
  assign storeAddrNotKnownFlags_12_2 = _T_16811 & entriesToCheck_12_2; // @[AxiLoadQueue.scala 163:19:@14151.4]
  assign storeAddrNotKnownFlags_12_3 = _T_16814 & entriesToCheck_12_3; // @[AxiLoadQueue.scala 163:19:@14153.4]
  assign storeAddrNotKnownFlags_12_4 = _T_16817 & entriesToCheck_12_4; // @[AxiLoadQueue.scala 163:19:@14155.4]
  assign storeAddrNotKnownFlags_12_5 = _T_16820 & entriesToCheck_12_5; // @[AxiLoadQueue.scala 163:19:@14157.4]
  assign storeAddrNotKnownFlags_12_6 = _T_16823 & entriesToCheck_12_6; // @[AxiLoadQueue.scala 163:19:@14159.4]
  assign storeAddrNotKnownFlags_12_7 = _T_16826 & entriesToCheck_12_7; // @[AxiLoadQueue.scala 163:19:@14161.4]
  assign storeAddrNotKnownFlags_12_8 = _T_16829 & entriesToCheck_12_8; // @[AxiLoadQueue.scala 163:19:@14163.4]
  assign storeAddrNotKnownFlags_12_9 = _T_16832 & entriesToCheck_12_9; // @[AxiLoadQueue.scala 163:19:@14165.4]
  assign storeAddrNotKnownFlags_12_10 = _T_16835 & entriesToCheck_12_10; // @[AxiLoadQueue.scala 163:19:@14167.4]
  assign storeAddrNotKnownFlags_12_11 = _T_16838 & entriesToCheck_12_11; // @[AxiLoadQueue.scala 163:19:@14169.4]
  assign storeAddrNotKnownFlags_12_12 = _T_16841 & entriesToCheck_12_12; // @[AxiLoadQueue.scala 163:19:@14171.4]
  assign storeAddrNotKnownFlags_12_13 = _T_16844 & entriesToCheck_12_13; // @[AxiLoadQueue.scala 163:19:@14173.4]
  assign storeAddrNotKnownFlags_12_14 = _T_16847 & entriesToCheck_12_14; // @[AxiLoadQueue.scala 163:19:@14175.4]
  assign storeAddrNotKnownFlags_12_15 = _T_16850 & entriesToCheck_12_15; // @[AxiLoadQueue.scala 163:19:@14177.4]
  assign storeAddrNotKnownFlags_13_0 = _T_16805 & entriesToCheck_13_0; // @[AxiLoadQueue.scala 163:19:@14195.4]
  assign storeAddrNotKnownFlags_13_1 = _T_16808 & entriesToCheck_13_1; // @[AxiLoadQueue.scala 163:19:@14197.4]
  assign storeAddrNotKnownFlags_13_2 = _T_16811 & entriesToCheck_13_2; // @[AxiLoadQueue.scala 163:19:@14199.4]
  assign storeAddrNotKnownFlags_13_3 = _T_16814 & entriesToCheck_13_3; // @[AxiLoadQueue.scala 163:19:@14201.4]
  assign storeAddrNotKnownFlags_13_4 = _T_16817 & entriesToCheck_13_4; // @[AxiLoadQueue.scala 163:19:@14203.4]
  assign storeAddrNotKnownFlags_13_5 = _T_16820 & entriesToCheck_13_5; // @[AxiLoadQueue.scala 163:19:@14205.4]
  assign storeAddrNotKnownFlags_13_6 = _T_16823 & entriesToCheck_13_6; // @[AxiLoadQueue.scala 163:19:@14207.4]
  assign storeAddrNotKnownFlags_13_7 = _T_16826 & entriesToCheck_13_7; // @[AxiLoadQueue.scala 163:19:@14209.4]
  assign storeAddrNotKnownFlags_13_8 = _T_16829 & entriesToCheck_13_8; // @[AxiLoadQueue.scala 163:19:@14211.4]
  assign storeAddrNotKnownFlags_13_9 = _T_16832 & entriesToCheck_13_9; // @[AxiLoadQueue.scala 163:19:@14213.4]
  assign storeAddrNotKnownFlags_13_10 = _T_16835 & entriesToCheck_13_10; // @[AxiLoadQueue.scala 163:19:@14215.4]
  assign storeAddrNotKnownFlags_13_11 = _T_16838 & entriesToCheck_13_11; // @[AxiLoadQueue.scala 163:19:@14217.4]
  assign storeAddrNotKnownFlags_13_12 = _T_16841 & entriesToCheck_13_12; // @[AxiLoadQueue.scala 163:19:@14219.4]
  assign storeAddrNotKnownFlags_13_13 = _T_16844 & entriesToCheck_13_13; // @[AxiLoadQueue.scala 163:19:@14221.4]
  assign storeAddrNotKnownFlags_13_14 = _T_16847 & entriesToCheck_13_14; // @[AxiLoadQueue.scala 163:19:@14223.4]
  assign storeAddrNotKnownFlags_13_15 = _T_16850 & entriesToCheck_13_15; // @[AxiLoadQueue.scala 163:19:@14225.4]
  assign storeAddrNotKnownFlags_14_0 = _T_16805 & entriesToCheck_14_0; // @[AxiLoadQueue.scala 163:19:@14243.4]
  assign storeAddrNotKnownFlags_14_1 = _T_16808 & entriesToCheck_14_1; // @[AxiLoadQueue.scala 163:19:@14245.4]
  assign storeAddrNotKnownFlags_14_2 = _T_16811 & entriesToCheck_14_2; // @[AxiLoadQueue.scala 163:19:@14247.4]
  assign storeAddrNotKnownFlags_14_3 = _T_16814 & entriesToCheck_14_3; // @[AxiLoadQueue.scala 163:19:@14249.4]
  assign storeAddrNotKnownFlags_14_4 = _T_16817 & entriesToCheck_14_4; // @[AxiLoadQueue.scala 163:19:@14251.4]
  assign storeAddrNotKnownFlags_14_5 = _T_16820 & entriesToCheck_14_5; // @[AxiLoadQueue.scala 163:19:@14253.4]
  assign storeAddrNotKnownFlags_14_6 = _T_16823 & entriesToCheck_14_6; // @[AxiLoadQueue.scala 163:19:@14255.4]
  assign storeAddrNotKnownFlags_14_7 = _T_16826 & entriesToCheck_14_7; // @[AxiLoadQueue.scala 163:19:@14257.4]
  assign storeAddrNotKnownFlags_14_8 = _T_16829 & entriesToCheck_14_8; // @[AxiLoadQueue.scala 163:19:@14259.4]
  assign storeAddrNotKnownFlags_14_9 = _T_16832 & entriesToCheck_14_9; // @[AxiLoadQueue.scala 163:19:@14261.4]
  assign storeAddrNotKnownFlags_14_10 = _T_16835 & entriesToCheck_14_10; // @[AxiLoadQueue.scala 163:19:@14263.4]
  assign storeAddrNotKnownFlags_14_11 = _T_16838 & entriesToCheck_14_11; // @[AxiLoadQueue.scala 163:19:@14265.4]
  assign storeAddrNotKnownFlags_14_12 = _T_16841 & entriesToCheck_14_12; // @[AxiLoadQueue.scala 163:19:@14267.4]
  assign storeAddrNotKnownFlags_14_13 = _T_16844 & entriesToCheck_14_13; // @[AxiLoadQueue.scala 163:19:@14269.4]
  assign storeAddrNotKnownFlags_14_14 = _T_16847 & entriesToCheck_14_14; // @[AxiLoadQueue.scala 163:19:@14271.4]
  assign storeAddrNotKnownFlags_14_15 = _T_16850 & entriesToCheck_14_15; // @[AxiLoadQueue.scala 163:19:@14273.4]
  assign storeAddrNotKnownFlags_15_0 = _T_16805 & entriesToCheck_15_0; // @[AxiLoadQueue.scala 163:19:@14291.4]
  assign storeAddrNotKnownFlags_15_1 = _T_16808 & entriesToCheck_15_1; // @[AxiLoadQueue.scala 163:19:@14293.4]
  assign storeAddrNotKnownFlags_15_2 = _T_16811 & entriesToCheck_15_2; // @[AxiLoadQueue.scala 163:19:@14295.4]
  assign storeAddrNotKnownFlags_15_3 = _T_16814 & entriesToCheck_15_3; // @[AxiLoadQueue.scala 163:19:@14297.4]
  assign storeAddrNotKnownFlags_15_4 = _T_16817 & entriesToCheck_15_4; // @[AxiLoadQueue.scala 163:19:@14299.4]
  assign storeAddrNotKnownFlags_15_5 = _T_16820 & entriesToCheck_15_5; // @[AxiLoadQueue.scala 163:19:@14301.4]
  assign storeAddrNotKnownFlags_15_6 = _T_16823 & entriesToCheck_15_6; // @[AxiLoadQueue.scala 163:19:@14303.4]
  assign storeAddrNotKnownFlags_15_7 = _T_16826 & entriesToCheck_15_7; // @[AxiLoadQueue.scala 163:19:@14305.4]
  assign storeAddrNotKnownFlags_15_8 = _T_16829 & entriesToCheck_15_8; // @[AxiLoadQueue.scala 163:19:@14307.4]
  assign storeAddrNotKnownFlags_15_9 = _T_16832 & entriesToCheck_15_9; // @[AxiLoadQueue.scala 163:19:@14309.4]
  assign storeAddrNotKnownFlags_15_10 = _T_16835 & entriesToCheck_15_10; // @[AxiLoadQueue.scala 163:19:@14311.4]
  assign storeAddrNotKnownFlags_15_11 = _T_16838 & entriesToCheck_15_11; // @[AxiLoadQueue.scala 163:19:@14313.4]
  assign storeAddrNotKnownFlags_15_12 = _T_16841 & entriesToCheck_15_12; // @[AxiLoadQueue.scala 163:19:@14315.4]
  assign storeAddrNotKnownFlags_15_13 = _T_16844 & entriesToCheck_15_13; // @[AxiLoadQueue.scala 163:19:@14317.4]
  assign storeAddrNotKnownFlags_15_14 = _T_16847 & entriesToCheck_15_14; // @[AxiLoadQueue.scala 163:19:@14319.4]
  assign storeAddrNotKnownFlags_15_15 = _T_16850 & entriesToCheck_15_15; // @[AxiLoadQueue.scala 163:19:@14321.4]
  assign _T_18008 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0}; // @[Mux.scala 19:72:@14652.4]
  assign _T_18015 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8}; // @[Mux.scala 19:72:@14659.4]
  assign _T_18016 = {conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,_T_18008}; // @[Mux.scala 19:72:@14660.4]
  assign _T_18018 = _T_2695 ? _T_18016 : 16'h0; // @[Mux.scala 19:72:@14661.4]
  assign _T_18025 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1}; // @[Mux.scala 19:72:@14668.4]
  assign _T_18032 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9}; // @[Mux.scala 19:72:@14675.4]
  assign _T_18033 = {conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,_T_18025}; // @[Mux.scala 19:72:@14676.4]
  assign _T_18035 = _T_2696 ? _T_18033 : 16'h0; // @[Mux.scala 19:72:@14677.4]
  assign _T_18042 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2}; // @[Mux.scala 19:72:@14684.4]
  assign _T_18049 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10}; // @[Mux.scala 19:72:@14691.4]
  assign _T_18050 = {conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,_T_18042}; // @[Mux.scala 19:72:@14692.4]
  assign _T_18052 = _T_2697 ? _T_18050 : 16'h0; // @[Mux.scala 19:72:@14693.4]
  assign _T_18059 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3}; // @[Mux.scala 19:72:@14700.4]
  assign _T_18066 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11}; // @[Mux.scala 19:72:@14707.4]
  assign _T_18067 = {conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,_T_18059}; // @[Mux.scala 19:72:@14708.4]
  assign _T_18069 = _T_2698 ? _T_18067 : 16'h0; // @[Mux.scala 19:72:@14709.4]
  assign _T_18076 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4}; // @[Mux.scala 19:72:@14716.4]
  assign _T_18083 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12}; // @[Mux.scala 19:72:@14723.4]
  assign _T_18084 = {conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,conflict_0_12,_T_18076}; // @[Mux.scala 19:72:@14724.4]
  assign _T_18086 = _T_2699 ? _T_18084 : 16'h0; // @[Mux.scala 19:72:@14725.4]
  assign _T_18093 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5}; // @[Mux.scala 19:72:@14732.4]
  assign _T_18100 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13}; // @[Mux.scala 19:72:@14739.4]
  assign _T_18101 = {conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,conflict_0_13,_T_18093}; // @[Mux.scala 19:72:@14740.4]
  assign _T_18103 = _T_2700 ? _T_18101 : 16'h0; // @[Mux.scala 19:72:@14741.4]
  assign _T_18110 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6}; // @[Mux.scala 19:72:@14748.4]
  assign _T_18117 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14}; // @[Mux.scala 19:72:@14755.4]
  assign _T_18118 = {conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,conflict_0_14,_T_18110}; // @[Mux.scala 19:72:@14756.4]
  assign _T_18120 = _T_2701 ? _T_18118 : 16'h0; // @[Mux.scala 19:72:@14757.4]
  assign _T_18127 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7}; // @[Mux.scala 19:72:@14764.4]
  assign _T_18134 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15}; // @[Mux.scala 19:72:@14771.4]
  assign _T_18135 = {conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,conflict_0_15,_T_18127}; // @[Mux.scala 19:72:@14772.4]
  assign _T_18137 = _T_2702 ? _T_18135 : 16'h0; // @[Mux.scala 19:72:@14773.4]
  assign _T_18152 = {conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,conflict_0_0,_T_18015}; // @[Mux.scala 19:72:@14788.4]
  assign _T_18154 = _T_2703 ? _T_18152 : 16'h0; // @[Mux.scala 19:72:@14789.4]
  assign _T_18169 = {conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,conflict_0_1,_T_18032}; // @[Mux.scala 19:72:@14804.4]
  assign _T_18171 = _T_2704 ? _T_18169 : 16'h0; // @[Mux.scala 19:72:@14805.4]
  assign _T_18186 = {conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,conflict_0_2,_T_18049}; // @[Mux.scala 19:72:@14820.4]
  assign _T_18188 = _T_2705 ? _T_18186 : 16'h0; // @[Mux.scala 19:72:@14821.4]
  assign _T_18203 = {conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,conflict_0_3,_T_18066}; // @[Mux.scala 19:72:@14836.4]
  assign _T_18205 = _T_2706 ? _T_18203 : 16'h0; // @[Mux.scala 19:72:@14837.4]
  assign _T_18220 = {conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,conflict_0_4,_T_18083}; // @[Mux.scala 19:72:@14852.4]
  assign _T_18222 = _T_2707 ? _T_18220 : 16'h0; // @[Mux.scala 19:72:@14853.4]
  assign _T_18237 = {conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,conflict_0_5,_T_18100}; // @[Mux.scala 19:72:@14868.4]
  assign _T_18239 = _T_2708 ? _T_18237 : 16'h0; // @[Mux.scala 19:72:@14869.4]
  assign _T_18254 = {conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,conflict_0_6,_T_18117}; // @[Mux.scala 19:72:@14884.4]
  assign _T_18256 = _T_2709 ? _T_18254 : 16'h0; // @[Mux.scala 19:72:@14885.4]
  assign _T_18271 = {conflict_0_14,conflict_0_13,conflict_0_12,conflict_0_11,conflict_0_10,conflict_0_9,conflict_0_8,conflict_0_7,_T_18134}; // @[Mux.scala 19:72:@14900.4]
  assign _T_18273 = _T_2710 ? _T_18271 : 16'h0; // @[Mux.scala 19:72:@14901.4]
  assign _T_18274 = _T_18018 | _T_18035; // @[Mux.scala 19:72:@14902.4]
  assign _T_18275 = _T_18274 | _T_18052; // @[Mux.scala 19:72:@14903.4]
  assign _T_18276 = _T_18275 | _T_18069; // @[Mux.scala 19:72:@14904.4]
  assign _T_18277 = _T_18276 | _T_18086; // @[Mux.scala 19:72:@14905.4]
  assign _T_18278 = _T_18277 | _T_18103; // @[Mux.scala 19:72:@14906.4]
  assign _T_18279 = _T_18278 | _T_18120; // @[Mux.scala 19:72:@14907.4]
  assign _T_18280 = _T_18279 | _T_18137; // @[Mux.scala 19:72:@14908.4]
  assign _T_18281 = _T_18280 | _T_18154; // @[Mux.scala 19:72:@14909.4]
  assign _T_18282 = _T_18281 | _T_18171; // @[Mux.scala 19:72:@14910.4]
  assign _T_18283 = _T_18282 | _T_18188; // @[Mux.scala 19:72:@14911.4]
  assign _T_18284 = _T_18283 | _T_18205; // @[Mux.scala 19:72:@14912.4]
  assign _T_18285 = _T_18284 | _T_18222; // @[Mux.scala 19:72:@14913.4]
  assign _T_18286 = _T_18285 | _T_18239; // @[Mux.scala 19:72:@14914.4]
  assign _T_18287 = _T_18286 | _T_18256; // @[Mux.scala 19:72:@14915.4]
  assign _T_18288 = _T_18287 | _T_18273; // @[Mux.scala 19:72:@14916.4]
  assign _T_18866 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0}; // @[Mux.scala 19:72:@15266.4]
  assign _T_18873 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8}; // @[Mux.scala 19:72:@15273.4]
  assign _T_18874 = {conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,_T_18866}; // @[Mux.scala 19:72:@15274.4]
  assign _T_18876 = _T_2695 ? _T_18874 : 16'h0; // @[Mux.scala 19:72:@15275.4]
  assign _T_18883 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1}; // @[Mux.scala 19:72:@15282.4]
  assign _T_18890 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9}; // @[Mux.scala 19:72:@15289.4]
  assign _T_18891 = {conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,_T_18883}; // @[Mux.scala 19:72:@15290.4]
  assign _T_18893 = _T_2696 ? _T_18891 : 16'h0; // @[Mux.scala 19:72:@15291.4]
  assign _T_18900 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2}; // @[Mux.scala 19:72:@15298.4]
  assign _T_18907 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10}; // @[Mux.scala 19:72:@15305.4]
  assign _T_18908 = {conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,_T_18900}; // @[Mux.scala 19:72:@15306.4]
  assign _T_18910 = _T_2697 ? _T_18908 : 16'h0; // @[Mux.scala 19:72:@15307.4]
  assign _T_18917 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3}; // @[Mux.scala 19:72:@15314.4]
  assign _T_18924 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11}; // @[Mux.scala 19:72:@15321.4]
  assign _T_18925 = {conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,_T_18917}; // @[Mux.scala 19:72:@15322.4]
  assign _T_18927 = _T_2698 ? _T_18925 : 16'h0; // @[Mux.scala 19:72:@15323.4]
  assign _T_18934 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4}; // @[Mux.scala 19:72:@15330.4]
  assign _T_18941 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12}; // @[Mux.scala 19:72:@15337.4]
  assign _T_18942 = {conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,conflict_1_12,_T_18934}; // @[Mux.scala 19:72:@15338.4]
  assign _T_18944 = _T_2699 ? _T_18942 : 16'h0; // @[Mux.scala 19:72:@15339.4]
  assign _T_18951 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5}; // @[Mux.scala 19:72:@15346.4]
  assign _T_18958 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13}; // @[Mux.scala 19:72:@15353.4]
  assign _T_18959 = {conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,conflict_1_13,_T_18951}; // @[Mux.scala 19:72:@15354.4]
  assign _T_18961 = _T_2700 ? _T_18959 : 16'h0; // @[Mux.scala 19:72:@15355.4]
  assign _T_18968 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6}; // @[Mux.scala 19:72:@15362.4]
  assign _T_18975 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14}; // @[Mux.scala 19:72:@15369.4]
  assign _T_18976 = {conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,conflict_1_14,_T_18968}; // @[Mux.scala 19:72:@15370.4]
  assign _T_18978 = _T_2701 ? _T_18976 : 16'h0; // @[Mux.scala 19:72:@15371.4]
  assign _T_18985 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7}; // @[Mux.scala 19:72:@15378.4]
  assign _T_18992 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15}; // @[Mux.scala 19:72:@15385.4]
  assign _T_18993 = {conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,conflict_1_15,_T_18985}; // @[Mux.scala 19:72:@15386.4]
  assign _T_18995 = _T_2702 ? _T_18993 : 16'h0; // @[Mux.scala 19:72:@15387.4]
  assign _T_19010 = {conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,conflict_1_0,_T_18873}; // @[Mux.scala 19:72:@15402.4]
  assign _T_19012 = _T_2703 ? _T_19010 : 16'h0; // @[Mux.scala 19:72:@15403.4]
  assign _T_19027 = {conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,conflict_1_1,_T_18890}; // @[Mux.scala 19:72:@15418.4]
  assign _T_19029 = _T_2704 ? _T_19027 : 16'h0; // @[Mux.scala 19:72:@15419.4]
  assign _T_19044 = {conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,conflict_1_2,_T_18907}; // @[Mux.scala 19:72:@15434.4]
  assign _T_19046 = _T_2705 ? _T_19044 : 16'h0; // @[Mux.scala 19:72:@15435.4]
  assign _T_19061 = {conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,conflict_1_3,_T_18924}; // @[Mux.scala 19:72:@15450.4]
  assign _T_19063 = _T_2706 ? _T_19061 : 16'h0; // @[Mux.scala 19:72:@15451.4]
  assign _T_19078 = {conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,conflict_1_4,_T_18941}; // @[Mux.scala 19:72:@15466.4]
  assign _T_19080 = _T_2707 ? _T_19078 : 16'h0; // @[Mux.scala 19:72:@15467.4]
  assign _T_19095 = {conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,conflict_1_5,_T_18958}; // @[Mux.scala 19:72:@15482.4]
  assign _T_19097 = _T_2708 ? _T_19095 : 16'h0; // @[Mux.scala 19:72:@15483.4]
  assign _T_19112 = {conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,conflict_1_6,_T_18975}; // @[Mux.scala 19:72:@15498.4]
  assign _T_19114 = _T_2709 ? _T_19112 : 16'h0; // @[Mux.scala 19:72:@15499.4]
  assign _T_19129 = {conflict_1_14,conflict_1_13,conflict_1_12,conflict_1_11,conflict_1_10,conflict_1_9,conflict_1_8,conflict_1_7,_T_18992}; // @[Mux.scala 19:72:@15514.4]
  assign _T_19131 = _T_2710 ? _T_19129 : 16'h0; // @[Mux.scala 19:72:@15515.4]
  assign _T_19132 = _T_18876 | _T_18893; // @[Mux.scala 19:72:@15516.4]
  assign _T_19133 = _T_19132 | _T_18910; // @[Mux.scala 19:72:@15517.4]
  assign _T_19134 = _T_19133 | _T_18927; // @[Mux.scala 19:72:@15518.4]
  assign _T_19135 = _T_19134 | _T_18944; // @[Mux.scala 19:72:@15519.4]
  assign _T_19136 = _T_19135 | _T_18961; // @[Mux.scala 19:72:@15520.4]
  assign _T_19137 = _T_19136 | _T_18978; // @[Mux.scala 19:72:@15521.4]
  assign _T_19138 = _T_19137 | _T_18995; // @[Mux.scala 19:72:@15522.4]
  assign _T_19139 = _T_19138 | _T_19012; // @[Mux.scala 19:72:@15523.4]
  assign _T_19140 = _T_19139 | _T_19029; // @[Mux.scala 19:72:@15524.4]
  assign _T_19141 = _T_19140 | _T_19046; // @[Mux.scala 19:72:@15525.4]
  assign _T_19142 = _T_19141 | _T_19063; // @[Mux.scala 19:72:@15526.4]
  assign _T_19143 = _T_19142 | _T_19080; // @[Mux.scala 19:72:@15527.4]
  assign _T_19144 = _T_19143 | _T_19097; // @[Mux.scala 19:72:@15528.4]
  assign _T_19145 = _T_19144 | _T_19114; // @[Mux.scala 19:72:@15529.4]
  assign _T_19146 = _T_19145 | _T_19131; // @[Mux.scala 19:72:@15530.4]
  assign _T_19724 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0}; // @[Mux.scala 19:72:@15880.4]
  assign _T_19731 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8}; // @[Mux.scala 19:72:@15887.4]
  assign _T_19732 = {conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,_T_19724}; // @[Mux.scala 19:72:@15888.4]
  assign _T_19734 = _T_2695 ? _T_19732 : 16'h0; // @[Mux.scala 19:72:@15889.4]
  assign _T_19741 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1}; // @[Mux.scala 19:72:@15896.4]
  assign _T_19748 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9}; // @[Mux.scala 19:72:@15903.4]
  assign _T_19749 = {conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,_T_19741}; // @[Mux.scala 19:72:@15904.4]
  assign _T_19751 = _T_2696 ? _T_19749 : 16'h0; // @[Mux.scala 19:72:@15905.4]
  assign _T_19758 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2}; // @[Mux.scala 19:72:@15912.4]
  assign _T_19765 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10}; // @[Mux.scala 19:72:@15919.4]
  assign _T_19766 = {conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,_T_19758}; // @[Mux.scala 19:72:@15920.4]
  assign _T_19768 = _T_2697 ? _T_19766 : 16'h0; // @[Mux.scala 19:72:@15921.4]
  assign _T_19775 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3}; // @[Mux.scala 19:72:@15928.4]
  assign _T_19782 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11}; // @[Mux.scala 19:72:@15935.4]
  assign _T_19783 = {conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,_T_19775}; // @[Mux.scala 19:72:@15936.4]
  assign _T_19785 = _T_2698 ? _T_19783 : 16'h0; // @[Mux.scala 19:72:@15937.4]
  assign _T_19792 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4}; // @[Mux.scala 19:72:@15944.4]
  assign _T_19799 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12}; // @[Mux.scala 19:72:@15951.4]
  assign _T_19800 = {conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,conflict_2_12,_T_19792}; // @[Mux.scala 19:72:@15952.4]
  assign _T_19802 = _T_2699 ? _T_19800 : 16'h0; // @[Mux.scala 19:72:@15953.4]
  assign _T_19809 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5}; // @[Mux.scala 19:72:@15960.4]
  assign _T_19816 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13}; // @[Mux.scala 19:72:@15967.4]
  assign _T_19817 = {conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,conflict_2_13,_T_19809}; // @[Mux.scala 19:72:@15968.4]
  assign _T_19819 = _T_2700 ? _T_19817 : 16'h0; // @[Mux.scala 19:72:@15969.4]
  assign _T_19826 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6}; // @[Mux.scala 19:72:@15976.4]
  assign _T_19833 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14}; // @[Mux.scala 19:72:@15983.4]
  assign _T_19834 = {conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,conflict_2_14,_T_19826}; // @[Mux.scala 19:72:@15984.4]
  assign _T_19836 = _T_2701 ? _T_19834 : 16'h0; // @[Mux.scala 19:72:@15985.4]
  assign _T_19843 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7}; // @[Mux.scala 19:72:@15992.4]
  assign _T_19850 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15}; // @[Mux.scala 19:72:@15999.4]
  assign _T_19851 = {conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,conflict_2_15,_T_19843}; // @[Mux.scala 19:72:@16000.4]
  assign _T_19853 = _T_2702 ? _T_19851 : 16'h0; // @[Mux.scala 19:72:@16001.4]
  assign _T_19868 = {conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,conflict_2_0,_T_19731}; // @[Mux.scala 19:72:@16016.4]
  assign _T_19870 = _T_2703 ? _T_19868 : 16'h0; // @[Mux.scala 19:72:@16017.4]
  assign _T_19885 = {conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,conflict_2_1,_T_19748}; // @[Mux.scala 19:72:@16032.4]
  assign _T_19887 = _T_2704 ? _T_19885 : 16'h0; // @[Mux.scala 19:72:@16033.4]
  assign _T_19902 = {conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,conflict_2_2,_T_19765}; // @[Mux.scala 19:72:@16048.4]
  assign _T_19904 = _T_2705 ? _T_19902 : 16'h0; // @[Mux.scala 19:72:@16049.4]
  assign _T_19919 = {conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,conflict_2_3,_T_19782}; // @[Mux.scala 19:72:@16064.4]
  assign _T_19921 = _T_2706 ? _T_19919 : 16'h0; // @[Mux.scala 19:72:@16065.4]
  assign _T_19936 = {conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,conflict_2_4,_T_19799}; // @[Mux.scala 19:72:@16080.4]
  assign _T_19938 = _T_2707 ? _T_19936 : 16'h0; // @[Mux.scala 19:72:@16081.4]
  assign _T_19953 = {conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,conflict_2_5,_T_19816}; // @[Mux.scala 19:72:@16096.4]
  assign _T_19955 = _T_2708 ? _T_19953 : 16'h0; // @[Mux.scala 19:72:@16097.4]
  assign _T_19970 = {conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,conflict_2_6,_T_19833}; // @[Mux.scala 19:72:@16112.4]
  assign _T_19972 = _T_2709 ? _T_19970 : 16'h0; // @[Mux.scala 19:72:@16113.4]
  assign _T_19987 = {conflict_2_14,conflict_2_13,conflict_2_12,conflict_2_11,conflict_2_10,conflict_2_9,conflict_2_8,conflict_2_7,_T_19850}; // @[Mux.scala 19:72:@16128.4]
  assign _T_19989 = _T_2710 ? _T_19987 : 16'h0; // @[Mux.scala 19:72:@16129.4]
  assign _T_19990 = _T_19734 | _T_19751; // @[Mux.scala 19:72:@16130.4]
  assign _T_19991 = _T_19990 | _T_19768; // @[Mux.scala 19:72:@16131.4]
  assign _T_19992 = _T_19991 | _T_19785; // @[Mux.scala 19:72:@16132.4]
  assign _T_19993 = _T_19992 | _T_19802; // @[Mux.scala 19:72:@16133.4]
  assign _T_19994 = _T_19993 | _T_19819; // @[Mux.scala 19:72:@16134.4]
  assign _T_19995 = _T_19994 | _T_19836; // @[Mux.scala 19:72:@16135.4]
  assign _T_19996 = _T_19995 | _T_19853; // @[Mux.scala 19:72:@16136.4]
  assign _T_19997 = _T_19996 | _T_19870; // @[Mux.scala 19:72:@16137.4]
  assign _T_19998 = _T_19997 | _T_19887; // @[Mux.scala 19:72:@16138.4]
  assign _T_19999 = _T_19998 | _T_19904; // @[Mux.scala 19:72:@16139.4]
  assign _T_20000 = _T_19999 | _T_19921; // @[Mux.scala 19:72:@16140.4]
  assign _T_20001 = _T_20000 | _T_19938; // @[Mux.scala 19:72:@16141.4]
  assign _T_20002 = _T_20001 | _T_19955; // @[Mux.scala 19:72:@16142.4]
  assign _T_20003 = _T_20002 | _T_19972; // @[Mux.scala 19:72:@16143.4]
  assign _T_20004 = _T_20003 | _T_19989; // @[Mux.scala 19:72:@16144.4]
  assign _T_20582 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0}; // @[Mux.scala 19:72:@16494.4]
  assign _T_20589 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8}; // @[Mux.scala 19:72:@16501.4]
  assign _T_20590 = {conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,_T_20582}; // @[Mux.scala 19:72:@16502.4]
  assign _T_20592 = _T_2695 ? _T_20590 : 16'h0; // @[Mux.scala 19:72:@16503.4]
  assign _T_20599 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1}; // @[Mux.scala 19:72:@16510.4]
  assign _T_20606 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9}; // @[Mux.scala 19:72:@16517.4]
  assign _T_20607 = {conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,_T_20599}; // @[Mux.scala 19:72:@16518.4]
  assign _T_20609 = _T_2696 ? _T_20607 : 16'h0; // @[Mux.scala 19:72:@16519.4]
  assign _T_20616 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2}; // @[Mux.scala 19:72:@16526.4]
  assign _T_20623 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10}; // @[Mux.scala 19:72:@16533.4]
  assign _T_20624 = {conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,_T_20616}; // @[Mux.scala 19:72:@16534.4]
  assign _T_20626 = _T_2697 ? _T_20624 : 16'h0; // @[Mux.scala 19:72:@16535.4]
  assign _T_20633 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3}; // @[Mux.scala 19:72:@16542.4]
  assign _T_20640 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11}; // @[Mux.scala 19:72:@16549.4]
  assign _T_20641 = {conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,_T_20633}; // @[Mux.scala 19:72:@16550.4]
  assign _T_20643 = _T_2698 ? _T_20641 : 16'h0; // @[Mux.scala 19:72:@16551.4]
  assign _T_20650 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4}; // @[Mux.scala 19:72:@16558.4]
  assign _T_20657 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12}; // @[Mux.scala 19:72:@16565.4]
  assign _T_20658 = {conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,conflict_3_12,_T_20650}; // @[Mux.scala 19:72:@16566.4]
  assign _T_20660 = _T_2699 ? _T_20658 : 16'h0; // @[Mux.scala 19:72:@16567.4]
  assign _T_20667 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5}; // @[Mux.scala 19:72:@16574.4]
  assign _T_20674 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13}; // @[Mux.scala 19:72:@16581.4]
  assign _T_20675 = {conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,conflict_3_13,_T_20667}; // @[Mux.scala 19:72:@16582.4]
  assign _T_20677 = _T_2700 ? _T_20675 : 16'h0; // @[Mux.scala 19:72:@16583.4]
  assign _T_20684 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6}; // @[Mux.scala 19:72:@16590.4]
  assign _T_20691 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14}; // @[Mux.scala 19:72:@16597.4]
  assign _T_20692 = {conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,conflict_3_14,_T_20684}; // @[Mux.scala 19:72:@16598.4]
  assign _T_20694 = _T_2701 ? _T_20692 : 16'h0; // @[Mux.scala 19:72:@16599.4]
  assign _T_20701 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7}; // @[Mux.scala 19:72:@16606.4]
  assign _T_20708 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15}; // @[Mux.scala 19:72:@16613.4]
  assign _T_20709 = {conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,conflict_3_15,_T_20701}; // @[Mux.scala 19:72:@16614.4]
  assign _T_20711 = _T_2702 ? _T_20709 : 16'h0; // @[Mux.scala 19:72:@16615.4]
  assign _T_20726 = {conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,conflict_3_0,_T_20589}; // @[Mux.scala 19:72:@16630.4]
  assign _T_20728 = _T_2703 ? _T_20726 : 16'h0; // @[Mux.scala 19:72:@16631.4]
  assign _T_20743 = {conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,conflict_3_1,_T_20606}; // @[Mux.scala 19:72:@16646.4]
  assign _T_20745 = _T_2704 ? _T_20743 : 16'h0; // @[Mux.scala 19:72:@16647.4]
  assign _T_20760 = {conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,conflict_3_2,_T_20623}; // @[Mux.scala 19:72:@16662.4]
  assign _T_20762 = _T_2705 ? _T_20760 : 16'h0; // @[Mux.scala 19:72:@16663.4]
  assign _T_20777 = {conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,conflict_3_3,_T_20640}; // @[Mux.scala 19:72:@16678.4]
  assign _T_20779 = _T_2706 ? _T_20777 : 16'h0; // @[Mux.scala 19:72:@16679.4]
  assign _T_20794 = {conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,conflict_3_4,_T_20657}; // @[Mux.scala 19:72:@16694.4]
  assign _T_20796 = _T_2707 ? _T_20794 : 16'h0; // @[Mux.scala 19:72:@16695.4]
  assign _T_20811 = {conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,conflict_3_5,_T_20674}; // @[Mux.scala 19:72:@16710.4]
  assign _T_20813 = _T_2708 ? _T_20811 : 16'h0; // @[Mux.scala 19:72:@16711.4]
  assign _T_20828 = {conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,conflict_3_6,_T_20691}; // @[Mux.scala 19:72:@16726.4]
  assign _T_20830 = _T_2709 ? _T_20828 : 16'h0; // @[Mux.scala 19:72:@16727.4]
  assign _T_20845 = {conflict_3_14,conflict_3_13,conflict_3_12,conflict_3_11,conflict_3_10,conflict_3_9,conflict_3_8,conflict_3_7,_T_20708}; // @[Mux.scala 19:72:@16742.4]
  assign _T_20847 = _T_2710 ? _T_20845 : 16'h0; // @[Mux.scala 19:72:@16743.4]
  assign _T_20848 = _T_20592 | _T_20609; // @[Mux.scala 19:72:@16744.4]
  assign _T_20849 = _T_20848 | _T_20626; // @[Mux.scala 19:72:@16745.4]
  assign _T_20850 = _T_20849 | _T_20643; // @[Mux.scala 19:72:@16746.4]
  assign _T_20851 = _T_20850 | _T_20660; // @[Mux.scala 19:72:@16747.4]
  assign _T_20852 = _T_20851 | _T_20677; // @[Mux.scala 19:72:@16748.4]
  assign _T_20853 = _T_20852 | _T_20694; // @[Mux.scala 19:72:@16749.4]
  assign _T_20854 = _T_20853 | _T_20711; // @[Mux.scala 19:72:@16750.4]
  assign _T_20855 = _T_20854 | _T_20728; // @[Mux.scala 19:72:@16751.4]
  assign _T_20856 = _T_20855 | _T_20745; // @[Mux.scala 19:72:@16752.4]
  assign _T_20857 = _T_20856 | _T_20762; // @[Mux.scala 19:72:@16753.4]
  assign _T_20858 = _T_20857 | _T_20779; // @[Mux.scala 19:72:@16754.4]
  assign _T_20859 = _T_20858 | _T_20796; // @[Mux.scala 19:72:@16755.4]
  assign _T_20860 = _T_20859 | _T_20813; // @[Mux.scala 19:72:@16756.4]
  assign _T_20861 = _T_20860 | _T_20830; // @[Mux.scala 19:72:@16757.4]
  assign _T_20862 = _T_20861 | _T_20847; // @[Mux.scala 19:72:@16758.4]
  assign _T_21440 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0}; // @[Mux.scala 19:72:@17108.4]
  assign _T_21447 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8}; // @[Mux.scala 19:72:@17115.4]
  assign _T_21448 = {conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,_T_21440}; // @[Mux.scala 19:72:@17116.4]
  assign _T_21450 = _T_2695 ? _T_21448 : 16'h0; // @[Mux.scala 19:72:@17117.4]
  assign _T_21457 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1}; // @[Mux.scala 19:72:@17124.4]
  assign _T_21464 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9}; // @[Mux.scala 19:72:@17131.4]
  assign _T_21465 = {conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,_T_21457}; // @[Mux.scala 19:72:@17132.4]
  assign _T_21467 = _T_2696 ? _T_21465 : 16'h0; // @[Mux.scala 19:72:@17133.4]
  assign _T_21474 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2}; // @[Mux.scala 19:72:@17140.4]
  assign _T_21481 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10}; // @[Mux.scala 19:72:@17147.4]
  assign _T_21482 = {conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,_T_21474}; // @[Mux.scala 19:72:@17148.4]
  assign _T_21484 = _T_2697 ? _T_21482 : 16'h0; // @[Mux.scala 19:72:@17149.4]
  assign _T_21491 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3}; // @[Mux.scala 19:72:@17156.4]
  assign _T_21498 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11}; // @[Mux.scala 19:72:@17163.4]
  assign _T_21499 = {conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,_T_21491}; // @[Mux.scala 19:72:@17164.4]
  assign _T_21501 = _T_2698 ? _T_21499 : 16'h0; // @[Mux.scala 19:72:@17165.4]
  assign _T_21508 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4}; // @[Mux.scala 19:72:@17172.4]
  assign _T_21515 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12}; // @[Mux.scala 19:72:@17179.4]
  assign _T_21516 = {conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,conflict_4_12,_T_21508}; // @[Mux.scala 19:72:@17180.4]
  assign _T_21518 = _T_2699 ? _T_21516 : 16'h0; // @[Mux.scala 19:72:@17181.4]
  assign _T_21525 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5}; // @[Mux.scala 19:72:@17188.4]
  assign _T_21532 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13}; // @[Mux.scala 19:72:@17195.4]
  assign _T_21533 = {conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,conflict_4_13,_T_21525}; // @[Mux.scala 19:72:@17196.4]
  assign _T_21535 = _T_2700 ? _T_21533 : 16'h0; // @[Mux.scala 19:72:@17197.4]
  assign _T_21542 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6}; // @[Mux.scala 19:72:@17204.4]
  assign _T_21549 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14}; // @[Mux.scala 19:72:@17211.4]
  assign _T_21550 = {conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,conflict_4_14,_T_21542}; // @[Mux.scala 19:72:@17212.4]
  assign _T_21552 = _T_2701 ? _T_21550 : 16'h0; // @[Mux.scala 19:72:@17213.4]
  assign _T_21559 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7}; // @[Mux.scala 19:72:@17220.4]
  assign _T_21566 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15}; // @[Mux.scala 19:72:@17227.4]
  assign _T_21567 = {conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,conflict_4_15,_T_21559}; // @[Mux.scala 19:72:@17228.4]
  assign _T_21569 = _T_2702 ? _T_21567 : 16'h0; // @[Mux.scala 19:72:@17229.4]
  assign _T_21584 = {conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,conflict_4_0,_T_21447}; // @[Mux.scala 19:72:@17244.4]
  assign _T_21586 = _T_2703 ? _T_21584 : 16'h0; // @[Mux.scala 19:72:@17245.4]
  assign _T_21601 = {conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,conflict_4_1,_T_21464}; // @[Mux.scala 19:72:@17260.4]
  assign _T_21603 = _T_2704 ? _T_21601 : 16'h0; // @[Mux.scala 19:72:@17261.4]
  assign _T_21618 = {conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,conflict_4_2,_T_21481}; // @[Mux.scala 19:72:@17276.4]
  assign _T_21620 = _T_2705 ? _T_21618 : 16'h0; // @[Mux.scala 19:72:@17277.4]
  assign _T_21635 = {conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,conflict_4_3,_T_21498}; // @[Mux.scala 19:72:@17292.4]
  assign _T_21637 = _T_2706 ? _T_21635 : 16'h0; // @[Mux.scala 19:72:@17293.4]
  assign _T_21652 = {conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,conflict_4_4,_T_21515}; // @[Mux.scala 19:72:@17308.4]
  assign _T_21654 = _T_2707 ? _T_21652 : 16'h0; // @[Mux.scala 19:72:@17309.4]
  assign _T_21669 = {conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,conflict_4_5,_T_21532}; // @[Mux.scala 19:72:@17324.4]
  assign _T_21671 = _T_2708 ? _T_21669 : 16'h0; // @[Mux.scala 19:72:@17325.4]
  assign _T_21686 = {conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,conflict_4_6,_T_21549}; // @[Mux.scala 19:72:@17340.4]
  assign _T_21688 = _T_2709 ? _T_21686 : 16'h0; // @[Mux.scala 19:72:@17341.4]
  assign _T_21703 = {conflict_4_14,conflict_4_13,conflict_4_12,conflict_4_11,conflict_4_10,conflict_4_9,conflict_4_8,conflict_4_7,_T_21566}; // @[Mux.scala 19:72:@17356.4]
  assign _T_21705 = _T_2710 ? _T_21703 : 16'h0; // @[Mux.scala 19:72:@17357.4]
  assign _T_21706 = _T_21450 | _T_21467; // @[Mux.scala 19:72:@17358.4]
  assign _T_21707 = _T_21706 | _T_21484; // @[Mux.scala 19:72:@17359.4]
  assign _T_21708 = _T_21707 | _T_21501; // @[Mux.scala 19:72:@17360.4]
  assign _T_21709 = _T_21708 | _T_21518; // @[Mux.scala 19:72:@17361.4]
  assign _T_21710 = _T_21709 | _T_21535; // @[Mux.scala 19:72:@17362.4]
  assign _T_21711 = _T_21710 | _T_21552; // @[Mux.scala 19:72:@17363.4]
  assign _T_21712 = _T_21711 | _T_21569; // @[Mux.scala 19:72:@17364.4]
  assign _T_21713 = _T_21712 | _T_21586; // @[Mux.scala 19:72:@17365.4]
  assign _T_21714 = _T_21713 | _T_21603; // @[Mux.scala 19:72:@17366.4]
  assign _T_21715 = _T_21714 | _T_21620; // @[Mux.scala 19:72:@17367.4]
  assign _T_21716 = _T_21715 | _T_21637; // @[Mux.scala 19:72:@17368.4]
  assign _T_21717 = _T_21716 | _T_21654; // @[Mux.scala 19:72:@17369.4]
  assign _T_21718 = _T_21717 | _T_21671; // @[Mux.scala 19:72:@17370.4]
  assign _T_21719 = _T_21718 | _T_21688; // @[Mux.scala 19:72:@17371.4]
  assign _T_21720 = _T_21719 | _T_21705; // @[Mux.scala 19:72:@17372.4]
  assign _T_22298 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0}; // @[Mux.scala 19:72:@17722.4]
  assign _T_22305 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8}; // @[Mux.scala 19:72:@17729.4]
  assign _T_22306 = {conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,_T_22298}; // @[Mux.scala 19:72:@17730.4]
  assign _T_22308 = _T_2695 ? _T_22306 : 16'h0; // @[Mux.scala 19:72:@17731.4]
  assign _T_22315 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1}; // @[Mux.scala 19:72:@17738.4]
  assign _T_22322 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9}; // @[Mux.scala 19:72:@17745.4]
  assign _T_22323 = {conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,_T_22315}; // @[Mux.scala 19:72:@17746.4]
  assign _T_22325 = _T_2696 ? _T_22323 : 16'h0; // @[Mux.scala 19:72:@17747.4]
  assign _T_22332 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2}; // @[Mux.scala 19:72:@17754.4]
  assign _T_22339 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10}; // @[Mux.scala 19:72:@17761.4]
  assign _T_22340 = {conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,_T_22332}; // @[Mux.scala 19:72:@17762.4]
  assign _T_22342 = _T_2697 ? _T_22340 : 16'h0; // @[Mux.scala 19:72:@17763.4]
  assign _T_22349 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3}; // @[Mux.scala 19:72:@17770.4]
  assign _T_22356 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11}; // @[Mux.scala 19:72:@17777.4]
  assign _T_22357 = {conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,_T_22349}; // @[Mux.scala 19:72:@17778.4]
  assign _T_22359 = _T_2698 ? _T_22357 : 16'h0; // @[Mux.scala 19:72:@17779.4]
  assign _T_22366 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4}; // @[Mux.scala 19:72:@17786.4]
  assign _T_22373 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12}; // @[Mux.scala 19:72:@17793.4]
  assign _T_22374 = {conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,conflict_5_12,_T_22366}; // @[Mux.scala 19:72:@17794.4]
  assign _T_22376 = _T_2699 ? _T_22374 : 16'h0; // @[Mux.scala 19:72:@17795.4]
  assign _T_22383 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5}; // @[Mux.scala 19:72:@17802.4]
  assign _T_22390 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13}; // @[Mux.scala 19:72:@17809.4]
  assign _T_22391 = {conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,conflict_5_13,_T_22383}; // @[Mux.scala 19:72:@17810.4]
  assign _T_22393 = _T_2700 ? _T_22391 : 16'h0; // @[Mux.scala 19:72:@17811.4]
  assign _T_22400 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6}; // @[Mux.scala 19:72:@17818.4]
  assign _T_22407 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14}; // @[Mux.scala 19:72:@17825.4]
  assign _T_22408 = {conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,conflict_5_14,_T_22400}; // @[Mux.scala 19:72:@17826.4]
  assign _T_22410 = _T_2701 ? _T_22408 : 16'h0; // @[Mux.scala 19:72:@17827.4]
  assign _T_22417 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7}; // @[Mux.scala 19:72:@17834.4]
  assign _T_22424 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15}; // @[Mux.scala 19:72:@17841.4]
  assign _T_22425 = {conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,conflict_5_15,_T_22417}; // @[Mux.scala 19:72:@17842.4]
  assign _T_22427 = _T_2702 ? _T_22425 : 16'h0; // @[Mux.scala 19:72:@17843.4]
  assign _T_22442 = {conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,conflict_5_0,_T_22305}; // @[Mux.scala 19:72:@17858.4]
  assign _T_22444 = _T_2703 ? _T_22442 : 16'h0; // @[Mux.scala 19:72:@17859.4]
  assign _T_22459 = {conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,conflict_5_1,_T_22322}; // @[Mux.scala 19:72:@17874.4]
  assign _T_22461 = _T_2704 ? _T_22459 : 16'h0; // @[Mux.scala 19:72:@17875.4]
  assign _T_22476 = {conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,conflict_5_2,_T_22339}; // @[Mux.scala 19:72:@17890.4]
  assign _T_22478 = _T_2705 ? _T_22476 : 16'h0; // @[Mux.scala 19:72:@17891.4]
  assign _T_22493 = {conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,conflict_5_3,_T_22356}; // @[Mux.scala 19:72:@17906.4]
  assign _T_22495 = _T_2706 ? _T_22493 : 16'h0; // @[Mux.scala 19:72:@17907.4]
  assign _T_22510 = {conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,conflict_5_4,_T_22373}; // @[Mux.scala 19:72:@17922.4]
  assign _T_22512 = _T_2707 ? _T_22510 : 16'h0; // @[Mux.scala 19:72:@17923.4]
  assign _T_22527 = {conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,conflict_5_5,_T_22390}; // @[Mux.scala 19:72:@17938.4]
  assign _T_22529 = _T_2708 ? _T_22527 : 16'h0; // @[Mux.scala 19:72:@17939.4]
  assign _T_22544 = {conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,conflict_5_6,_T_22407}; // @[Mux.scala 19:72:@17954.4]
  assign _T_22546 = _T_2709 ? _T_22544 : 16'h0; // @[Mux.scala 19:72:@17955.4]
  assign _T_22561 = {conflict_5_14,conflict_5_13,conflict_5_12,conflict_5_11,conflict_5_10,conflict_5_9,conflict_5_8,conflict_5_7,_T_22424}; // @[Mux.scala 19:72:@17970.4]
  assign _T_22563 = _T_2710 ? _T_22561 : 16'h0; // @[Mux.scala 19:72:@17971.4]
  assign _T_22564 = _T_22308 | _T_22325; // @[Mux.scala 19:72:@17972.4]
  assign _T_22565 = _T_22564 | _T_22342; // @[Mux.scala 19:72:@17973.4]
  assign _T_22566 = _T_22565 | _T_22359; // @[Mux.scala 19:72:@17974.4]
  assign _T_22567 = _T_22566 | _T_22376; // @[Mux.scala 19:72:@17975.4]
  assign _T_22568 = _T_22567 | _T_22393; // @[Mux.scala 19:72:@17976.4]
  assign _T_22569 = _T_22568 | _T_22410; // @[Mux.scala 19:72:@17977.4]
  assign _T_22570 = _T_22569 | _T_22427; // @[Mux.scala 19:72:@17978.4]
  assign _T_22571 = _T_22570 | _T_22444; // @[Mux.scala 19:72:@17979.4]
  assign _T_22572 = _T_22571 | _T_22461; // @[Mux.scala 19:72:@17980.4]
  assign _T_22573 = _T_22572 | _T_22478; // @[Mux.scala 19:72:@17981.4]
  assign _T_22574 = _T_22573 | _T_22495; // @[Mux.scala 19:72:@17982.4]
  assign _T_22575 = _T_22574 | _T_22512; // @[Mux.scala 19:72:@17983.4]
  assign _T_22576 = _T_22575 | _T_22529; // @[Mux.scala 19:72:@17984.4]
  assign _T_22577 = _T_22576 | _T_22546; // @[Mux.scala 19:72:@17985.4]
  assign _T_22578 = _T_22577 | _T_22563; // @[Mux.scala 19:72:@17986.4]
  assign _T_23156 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0}; // @[Mux.scala 19:72:@18336.4]
  assign _T_23163 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8}; // @[Mux.scala 19:72:@18343.4]
  assign _T_23164 = {conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,_T_23156}; // @[Mux.scala 19:72:@18344.4]
  assign _T_23166 = _T_2695 ? _T_23164 : 16'h0; // @[Mux.scala 19:72:@18345.4]
  assign _T_23173 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1}; // @[Mux.scala 19:72:@18352.4]
  assign _T_23180 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9}; // @[Mux.scala 19:72:@18359.4]
  assign _T_23181 = {conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,_T_23173}; // @[Mux.scala 19:72:@18360.4]
  assign _T_23183 = _T_2696 ? _T_23181 : 16'h0; // @[Mux.scala 19:72:@18361.4]
  assign _T_23190 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2}; // @[Mux.scala 19:72:@18368.4]
  assign _T_23197 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10}; // @[Mux.scala 19:72:@18375.4]
  assign _T_23198 = {conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,_T_23190}; // @[Mux.scala 19:72:@18376.4]
  assign _T_23200 = _T_2697 ? _T_23198 : 16'h0; // @[Mux.scala 19:72:@18377.4]
  assign _T_23207 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3}; // @[Mux.scala 19:72:@18384.4]
  assign _T_23214 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11}; // @[Mux.scala 19:72:@18391.4]
  assign _T_23215 = {conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,_T_23207}; // @[Mux.scala 19:72:@18392.4]
  assign _T_23217 = _T_2698 ? _T_23215 : 16'h0; // @[Mux.scala 19:72:@18393.4]
  assign _T_23224 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4}; // @[Mux.scala 19:72:@18400.4]
  assign _T_23231 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12}; // @[Mux.scala 19:72:@18407.4]
  assign _T_23232 = {conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,conflict_6_12,_T_23224}; // @[Mux.scala 19:72:@18408.4]
  assign _T_23234 = _T_2699 ? _T_23232 : 16'h0; // @[Mux.scala 19:72:@18409.4]
  assign _T_23241 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5}; // @[Mux.scala 19:72:@18416.4]
  assign _T_23248 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13}; // @[Mux.scala 19:72:@18423.4]
  assign _T_23249 = {conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,conflict_6_13,_T_23241}; // @[Mux.scala 19:72:@18424.4]
  assign _T_23251 = _T_2700 ? _T_23249 : 16'h0; // @[Mux.scala 19:72:@18425.4]
  assign _T_23258 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6}; // @[Mux.scala 19:72:@18432.4]
  assign _T_23265 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14}; // @[Mux.scala 19:72:@18439.4]
  assign _T_23266 = {conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,conflict_6_14,_T_23258}; // @[Mux.scala 19:72:@18440.4]
  assign _T_23268 = _T_2701 ? _T_23266 : 16'h0; // @[Mux.scala 19:72:@18441.4]
  assign _T_23275 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7}; // @[Mux.scala 19:72:@18448.4]
  assign _T_23282 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15}; // @[Mux.scala 19:72:@18455.4]
  assign _T_23283 = {conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,conflict_6_15,_T_23275}; // @[Mux.scala 19:72:@18456.4]
  assign _T_23285 = _T_2702 ? _T_23283 : 16'h0; // @[Mux.scala 19:72:@18457.4]
  assign _T_23300 = {conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,conflict_6_0,_T_23163}; // @[Mux.scala 19:72:@18472.4]
  assign _T_23302 = _T_2703 ? _T_23300 : 16'h0; // @[Mux.scala 19:72:@18473.4]
  assign _T_23317 = {conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,conflict_6_1,_T_23180}; // @[Mux.scala 19:72:@18488.4]
  assign _T_23319 = _T_2704 ? _T_23317 : 16'h0; // @[Mux.scala 19:72:@18489.4]
  assign _T_23334 = {conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,conflict_6_2,_T_23197}; // @[Mux.scala 19:72:@18504.4]
  assign _T_23336 = _T_2705 ? _T_23334 : 16'h0; // @[Mux.scala 19:72:@18505.4]
  assign _T_23351 = {conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,conflict_6_3,_T_23214}; // @[Mux.scala 19:72:@18520.4]
  assign _T_23353 = _T_2706 ? _T_23351 : 16'h0; // @[Mux.scala 19:72:@18521.4]
  assign _T_23368 = {conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,conflict_6_4,_T_23231}; // @[Mux.scala 19:72:@18536.4]
  assign _T_23370 = _T_2707 ? _T_23368 : 16'h0; // @[Mux.scala 19:72:@18537.4]
  assign _T_23385 = {conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,conflict_6_5,_T_23248}; // @[Mux.scala 19:72:@18552.4]
  assign _T_23387 = _T_2708 ? _T_23385 : 16'h0; // @[Mux.scala 19:72:@18553.4]
  assign _T_23402 = {conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,conflict_6_6,_T_23265}; // @[Mux.scala 19:72:@18568.4]
  assign _T_23404 = _T_2709 ? _T_23402 : 16'h0; // @[Mux.scala 19:72:@18569.4]
  assign _T_23419 = {conflict_6_14,conflict_6_13,conflict_6_12,conflict_6_11,conflict_6_10,conflict_6_9,conflict_6_8,conflict_6_7,_T_23282}; // @[Mux.scala 19:72:@18584.4]
  assign _T_23421 = _T_2710 ? _T_23419 : 16'h0; // @[Mux.scala 19:72:@18585.4]
  assign _T_23422 = _T_23166 | _T_23183; // @[Mux.scala 19:72:@18586.4]
  assign _T_23423 = _T_23422 | _T_23200; // @[Mux.scala 19:72:@18587.4]
  assign _T_23424 = _T_23423 | _T_23217; // @[Mux.scala 19:72:@18588.4]
  assign _T_23425 = _T_23424 | _T_23234; // @[Mux.scala 19:72:@18589.4]
  assign _T_23426 = _T_23425 | _T_23251; // @[Mux.scala 19:72:@18590.4]
  assign _T_23427 = _T_23426 | _T_23268; // @[Mux.scala 19:72:@18591.4]
  assign _T_23428 = _T_23427 | _T_23285; // @[Mux.scala 19:72:@18592.4]
  assign _T_23429 = _T_23428 | _T_23302; // @[Mux.scala 19:72:@18593.4]
  assign _T_23430 = _T_23429 | _T_23319; // @[Mux.scala 19:72:@18594.4]
  assign _T_23431 = _T_23430 | _T_23336; // @[Mux.scala 19:72:@18595.4]
  assign _T_23432 = _T_23431 | _T_23353; // @[Mux.scala 19:72:@18596.4]
  assign _T_23433 = _T_23432 | _T_23370; // @[Mux.scala 19:72:@18597.4]
  assign _T_23434 = _T_23433 | _T_23387; // @[Mux.scala 19:72:@18598.4]
  assign _T_23435 = _T_23434 | _T_23404; // @[Mux.scala 19:72:@18599.4]
  assign _T_23436 = _T_23435 | _T_23421; // @[Mux.scala 19:72:@18600.4]
  assign _T_24014 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0}; // @[Mux.scala 19:72:@18950.4]
  assign _T_24021 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8}; // @[Mux.scala 19:72:@18957.4]
  assign _T_24022 = {conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,_T_24014}; // @[Mux.scala 19:72:@18958.4]
  assign _T_24024 = _T_2695 ? _T_24022 : 16'h0; // @[Mux.scala 19:72:@18959.4]
  assign _T_24031 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1}; // @[Mux.scala 19:72:@18966.4]
  assign _T_24038 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9}; // @[Mux.scala 19:72:@18973.4]
  assign _T_24039 = {conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,_T_24031}; // @[Mux.scala 19:72:@18974.4]
  assign _T_24041 = _T_2696 ? _T_24039 : 16'h0; // @[Mux.scala 19:72:@18975.4]
  assign _T_24048 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2}; // @[Mux.scala 19:72:@18982.4]
  assign _T_24055 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10}; // @[Mux.scala 19:72:@18989.4]
  assign _T_24056 = {conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,_T_24048}; // @[Mux.scala 19:72:@18990.4]
  assign _T_24058 = _T_2697 ? _T_24056 : 16'h0; // @[Mux.scala 19:72:@18991.4]
  assign _T_24065 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3}; // @[Mux.scala 19:72:@18998.4]
  assign _T_24072 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11}; // @[Mux.scala 19:72:@19005.4]
  assign _T_24073 = {conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,_T_24065}; // @[Mux.scala 19:72:@19006.4]
  assign _T_24075 = _T_2698 ? _T_24073 : 16'h0; // @[Mux.scala 19:72:@19007.4]
  assign _T_24082 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4}; // @[Mux.scala 19:72:@19014.4]
  assign _T_24089 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12}; // @[Mux.scala 19:72:@19021.4]
  assign _T_24090 = {conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,conflict_7_12,_T_24082}; // @[Mux.scala 19:72:@19022.4]
  assign _T_24092 = _T_2699 ? _T_24090 : 16'h0; // @[Mux.scala 19:72:@19023.4]
  assign _T_24099 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5}; // @[Mux.scala 19:72:@19030.4]
  assign _T_24106 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13}; // @[Mux.scala 19:72:@19037.4]
  assign _T_24107 = {conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,conflict_7_13,_T_24099}; // @[Mux.scala 19:72:@19038.4]
  assign _T_24109 = _T_2700 ? _T_24107 : 16'h0; // @[Mux.scala 19:72:@19039.4]
  assign _T_24116 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6}; // @[Mux.scala 19:72:@19046.4]
  assign _T_24123 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14}; // @[Mux.scala 19:72:@19053.4]
  assign _T_24124 = {conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,conflict_7_14,_T_24116}; // @[Mux.scala 19:72:@19054.4]
  assign _T_24126 = _T_2701 ? _T_24124 : 16'h0; // @[Mux.scala 19:72:@19055.4]
  assign _T_24133 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7}; // @[Mux.scala 19:72:@19062.4]
  assign _T_24140 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15}; // @[Mux.scala 19:72:@19069.4]
  assign _T_24141 = {conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,conflict_7_15,_T_24133}; // @[Mux.scala 19:72:@19070.4]
  assign _T_24143 = _T_2702 ? _T_24141 : 16'h0; // @[Mux.scala 19:72:@19071.4]
  assign _T_24158 = {conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,conflict_7_0,_T_24021}; // @[Mux.scala 19:72:@19086.4]
  assign _T_24160 = _T_2703 ? _T_24158 : 16'h0; // @[Mux.scala 19:72:@19087.4]
  assign _T_24175 = {conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,conflict_7_1,_T_24038}; // @[Mux.scala 19:72:@19102.4]
  assign _T_24177 = _T_2704 ? _T_24175 : 16'h0; // @[Mux.scala 19:72:@19103.4]
  assign _T_24192 = {conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,conflict_7_2,_T_24055}; // @[Mux.scala 19:72:@19118.4]
  assign _T_24194 = _T_2705 ? _T_24192 : 16'h0; // @[Mux.scala 19:72:@19119.4]
  assign _T_24209 = {conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,conflict_7_3,_T_24072}; // @[Mux.scala 19:72:@19134.4]
  assign _T_24211 = _T_2706 ? _T_24209 : 16'h0; // @[Mux.scala 19:72:@19135.4]
  assign _T_24226 = {conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,conflict_7_4,_T_24089}; // @[Mux.scala 19:72:@19150.4]
  assign _T_24228 = _T_2707 ? _T_24226 : 16'h0; // @[Mux.scala 19:72:@19151.4]
  assign _T_24243 = {conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,conflict_7_5,_T_24106}; // @[Mux.scala 19:72:@19166.4]
  assign _T_24245 = _T_2708 ? _T_24243 : 16'h0; // @[Mux.scala 19:72:@19167.4]
  assign _T_24260 = {conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,conflict_7_6,_T_24123}; // @[Mux.scala 19:72:@19182.4]
  assign _T_24262 = _T_2709 ? _T_24260 : 16'h0; // @[Mux.scala 19:72:@19183.4]
  assign _T_24277 = {conflict_7_14,conflict_7_13,conflict_7_12,conflict_7_11,conflict_7_10,conflict_7_9,conflict_7_8,conflict_7_7,_T_24140}; // @[Mux.scala 19:72:@19198.4]
  assign _T_24279 = _T_2710 ? _T_24277 : 16'h0; // @[Mux.scala 19:72:@19199.4]
  assign _T_24280 = _T_24024 | _T_24041; // @[Mux.scala 19:72:@19200.4]
  assign _T_24281 = _T_24280 | _T_24058; // @[Mux.scala 19:72:@19201.4]
  assign _T_24282 = _T_24281 | _T_24075; // @[Mux.scala 19:72:@19202.4]
  assign _T_24283 = _T_24282 | _T_24092; // @[Mux.scala 19:72:@19203.4]
  assign _T_24284 = _T_24283 | _T_24109; // @[Mux.scala 19:72:@19204.4]
  assign _T_24285 = _T_24284 | _T_24126; // @[Mux.scala 19:72:@19205.4]
  assign _T_24286 = _T_24285 | _T_24143; // @[Mux.scala 19:72:@19206.4]
  assign _T_24287 = _T_24286 | _T_24160; // @[Mux.scala 19:72:@19207.4]
  assign _T_24288 = _T_24287 | _T_24177; // @[Mux.scala 19:72:@19208.4]
  assign _T_24289 = _T_24288 | _T_24194; // @[Mux.scala 19:72:@19209.4]
  assign _T_24290 = _T_24289 | _T_24211; // @[Mux.scala 19:72:@19210.4]
  assign _T_24291 = _T_24290 | _T_24228; // @[Mux.scala 19:72:@19211.4]
  assign _T_24292 = _T_24291 | _T_24245; // @[Mux.scala 19:72:@19212.4]
  assign _T_24293 = _T_24292 | _T_24262; // @[Mux.scala 19:72:@19213.4]
  assign _T_24294 = _T_24293 | _T_24279; // @[Mux.scala 19:72:@19214.4]
  assign _T_24872 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0}; // @[Mux.scala 19:72:@19564.4]
  assign _T_24879 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8}; // @[Mux.scala 19:72:@19571.4]
  assign _T_24880 = {conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,_T_24872}; // @[Mux.scala 19:72:@19572.4]
  assign _T_24882 = _T_2695 ? _T_24880 : 16'h0; // @[Mux.scala 19:72:@19573.4]
  assign _T_24889 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1}; // @[Mux.scala 19:72:@19580.4]
  assign _T_24896 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9}; // @[Mux.scala 19:72:@19587.4]
  assign _T_24897 = {conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,_T_24889}; // @[Mux.scala 19:72:@19588.4]
  assign _T_24899 = _T_2696 ? _T_24897 : 16'h0; // @[Mux.scala 19:72:@19589.4]
  assign _T_24906 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2}; // @[Mux.scala 19:72:@19596.4]
  assign _T_24913 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10}; // @[Mux.scala 19:72:@19603.4]
  assign _T_24914 = {conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,_T_24906}; // @[Mux.scala 19:72:@19604.4]
  assign _T_24916 = _T_2697 ? _T_24914 : 16'h0; // @[Mux.scala 19:72:@19605.4]
  assign _T_24923 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3}; // @[Mux.scala 19:72:@19612.4]
  assign _T_24930 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11}; // @[Mux.scala 19:72:@19619.4]
  assign _T_24931 = {conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,_T_24923}; // @[Mux.scala 19:72:@19620.4]
  assign _T_24933 = _T_2698 ? _T_24931 : 16'h0; // @[Mux.scala 19:72:@19621.4]
  assign _T_24940 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4}; // @[Mux.scala 19:72:@19628.4]
  assign _T_24947 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12}; // @[Mux.scala 19:72:@19635.4]
  assign _T_24948 = {conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,conflict_8_12,_T_24940}; // @[Mux.scala 19:72:@19636.4]
  assign _T_24950 = _T_2699 ? _T_24948 : 16'h0; // @[Mux.scala 19:72:@19637.4]
  assign _T_24957 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5}; // @[Mux.scala 19:72:@19644.4]
  assign _T_24964 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13}; // @[Mux.scala 19:72:@19651.4]
  assign _T_24965 = {conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,conflict_8_13,_T_24957}; // @[Mux.scala 19:72:@19652.4]
  assign _T_24967 = _T_2700 ? _T_24965 : 16'h0; // @[Mux.scala 19:72:@19653.4]
  assign _T_24974 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6}; // @[Mux.scala 19:72:@19660.4]
  assign _T_24981 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14}; // @[Mux.scala 19:72:@19667.4]
  assign _T_24982 = {conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,conflict_8_14,_T_24974}; // @[Mux.scala 19:72:@19668.4]
  assign _T_24984 = _T_2701 ? _T_24982 : 16'h0; // @[Mux.scala 19:72:@19669.4]
  assign _T_24991 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7}; // @[Mux.scala 19:72:@19676.4]
  assign _T_24998 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15}; // @[Mux.scala 19:72:@19683.4]
  assign _T_24999 = {conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,conflict_8_15,_T_24991}; // @[Mux.scala 19:72:@19684.4]
  assign _T_25001 = _T_2702 ? _T_24999 : 16'h0; // @[Mux.scala 19:72:@19685.4]
  assign _T_25016 = {conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,conflict_8_0,_T_24879}; // @[Mux.scala 19:72:@19700.4]
  assign _T_25018 = _T_2703 ? _T_25016 : 16'h0; // @[Mux.scala 19:72:@19701.4]
  assign _T_25033 = {conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,conflict_8_1,_T_24896}; // @[Mux.scala 19:72:@19716.4]
  assign _T_25035 = _T_2704 ? _T_25033 : 16'h0; // @[Mux.scala 19:72:@19717.4]
  assign _T_25050 = {conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,conflict_8_2,_T_24913}; // @[Mux.scala 19:72:@19732.4]
  assign _T_25052 = _T_2705 ? _T_25050 : 16'h0; // @[Mux.scala 19:72:@19733.4]
  assign _T_25067 = {conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,conflict_8_3,_T_24930}; // @[Mux.scala 19:72:@19748.4]
  assign _T_25069 = _T_2706 ? _T_25067 : 16'h0; // @[Mux.scala 19:72:@19749.4]
  assign _T_25084 = {conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,conflict_8_4,_T_24947}; // @[Mux.scala 19:72:@19764.4]
  assign _T_25086 = _T_2707 ? _T_25084 : 16'h0; // @[Mux.scala 19:72:@19765.4]
  assign _T_25101 = {conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,conflict_8_5,_T_24964}; // @[Mux.scala 19:72:@19780.4]
  assign _T_25103 = _T_2708 ? _T_25101 : 16'h0; // @[Mux.scala 19:72:@19781.4]
  assign _T_25118 = {conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,conflict_8_6,_T_24981}; // @[Mux.scala 19:72:@19796.4]
  assign _T_25120 = _T_2709 ? _T_25118 : 16'h0; // @[Mux.scala 19:72:@19797.4]
  assign _T_25135 = {conflict_8_14,conflict_8_13,conflict_8_12,conflict_8_11,conflict_8_10,conflict_8_9,conflict_8_8,conflict_8_7,_T_24998}; // @[Mux.scala 19:72:@19812.4]
  assign _T_25137 = _T_2710 ? _T_25135 : 16'h0; // @[Mux.scala 19:72:@19813.4]
  assign _T_25138 = _T_24882 | _T_24899; // @[Mux.scala 19:72:@19814.4]
  assign _T_25139 = _T_25138 | _T_24916; // @[Mux.scala 19:72:@19815.4]
  assign _T_25140 = _T_25139 | _T_24933; // @[Mux.scala 19:72:@19816.4]
  assign _T_25141 = _T_25140 | _T_24950; // @[Mux.scala 19:72:@19817.4]
  assign _T_25142 = _T_25141 | _T_24967; // @[Mux.scala 19:72:@19818.4]
  assign _T_25143 = _T_25142 | _T_24984; // @[Mux.scala 19:72:@19819.4]
  assign _T_25144 = _T_25143 | _T_25001; // @[Mux.scala 19:72:@19820.4]
  assign _T_25145 = _T_25144 | _T_25018; // @[Mux.scala 19:72:@19821.4]
  assign _T_25146 = _T_25145 | _T_25035; // @[Mux.scala 19:72:@19822.4]
  assign _T_25147 = _T_25146 | _T_25052; // @[Mux.scala 19:72:@19823.4]
  assign _T_25148 = _T_25147 | _T_25069; // @[Mux.scala 19:72:@19824.4]
  assign _T_25149 = _T_25148 | _T_25086; // @[Mux.scala 19:72:@19825.4]
  assign _T_25150 = _T_25149 | _T_25103; // @[Mux.scala 19:72:@19826.4]
  assign _T_25151 = _T_25150 | _T_25120; // @[Mux.scala 19:72:@19827.4]
  assign _T_25152 = _T_25151 | _T_25137; // @[Mux.scala 19:72:@19828.4]
  assign _T_25730 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0}; // @[Mux.scala 19:72:@20178.4]
  assign _T_25737 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8}; // @[Mux.scala 19:72:@20185.4]
  assign _T_25738 = {conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,_T_25730}; // @[Mux.scala 19:72:@20186.4]
  assign _T_25740 = _T_2695 ? _T_25738 : 16'h0; // @[Mux.scala 19:72:@20187.4]
  assign _T_25747 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1}; // @[Mux.scala 19:72:@20194.4]
  assign _T_25754 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9}; // @[Mux.scala 19:72:@20201.4]
  assign _T_25755 = {conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,_T_25747}; // @[Mux.scala 19:72:@20202.4]
  assign _T_25757 = _T_2696 ? _T_25755 : 16'h0; // @[Mux.scala 19:72:@20203.4]
  assign _T_25764 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2}; // @[Mux.scala 19:72:@20210.4]
  assign _T_25771 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10}; // @[Mux.scala 19:72:@20217.4]
  assign _T_25772 = {conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,_T_25764}; // @[Mux.scala 19:72:@20218.4]
  assign _T_25774 = _T_2697 ? _T_25772 : 16'h0; // @[Mux.scala 19:72:@20219.4]
  assign _T_25781 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3}; // @[Mux.scala 19:72:@20226.4]
  assign _T_25788 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11}; // @[Mux.scala 19:72:@20233.4]
  assign _T_25789 = {conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,_T_25781}; // @[Mux.scala 19:72:@20234.4]
  assign _T_25791 = _T_2698 ? _T_25789 : 16'h0; // @[Mux.scala 19:72:@20235.4]
  assign _T_25798 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4}; // @[Mux.scala 19:72:@20242.4]
  assign _T_25805 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12}; // @[Mux.scala 19:72:@20249.4]
  assign _T_25806 = {conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,conflict_9_12,_T_25798}; // @[Mux.scala 19:72:@20250.4]
  assign _T_25808 = _T_2699 ? _T_25806 : 16'h0; // @[Mux.scala 19:72:@20251.4]
  assign _T_25815 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5}; // @[Mux.scala 19:72:@20258.4]
  assign _T_25822 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13}; // @[Mux.scala 19:72:@20265.4]
  assign _T_25823 = {conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,conflict_9_13,_T_25815}; // @[Mux.scala 19:72:@20266.4]
  assign _T_25825 = _T_2700 ? _T_25823 : 16'h0; // @[Mux.scala 19:72:@20267.4]
  assign _T_25832 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6}; // @[Mux.scala 19:72:@20274.4]
  assign _T_25839 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14}; // @[Mux.scala 19:72:@20281.4]
  assign _T_25840 = {conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,conflict_9_14,_T_25832}; // @[Mux.scala 19:72:@20282.4]
  assign _T_25842 = _T_2701 ? _T_25840 : 16'h0; // @[Mux.scala 19:72:@20283.4]
  assign _T_25849 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7}; // @[Mux.scala 19:72:@20290.4]
  assign _T_25856 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15}; // @[Mux.scala 19:72:@20297.4]
  assign _T_25857 = {conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,conflict_9_15,_T_25849}; // @[Mux.scala 19:72:@20298.4]
  assign _T_25859 = _T_2702 ? _T_25857 : 16'h0; // @[Mux.scala 19:72:@20299.4]
  assign _T_25874 = {conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,conflict_9_0,_T_25737}; // @[Mux.scala 19:72:@20314.4]
  assign _T_25876 = _T_2703 ? _T_25874 : 16'h0; // @[Mux.scala 19:72:@20315.4]
  assign _T_25891 = {conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,conflict_9_1,_T_25754}; // @[Mux.scala 19:72:@20330.4]
  assign _T_25893 = _T_2704 ? _T_25891 : 16'h0; // @[Mux.scala 19:72:@20331.4]
  assign _T_25908 = {conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,conflict_9_2,_T_25771}; // @[Mux.scala 19:72:@20346.4]
  assign _T_25910 = _T_2705 ? _T_25908 : 16'h0; // @[Mux.scala 19:72:@20347.4]
  assign _T_25925 = {conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,conflict_9_3,_T_25788}; // @[Mux.scala 19:72:@20362.4]
  assign _T_25927 = _T_2706 ? _T_25925 : 16'h0; // @[Mux.scala 19:72:@20363.4]
  assign _T_25942 = {conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,conflict_9_4,_T_25805}; // @[Mux.scala 19:72:@20378.4]
  assign _T_25944 = _T_2707 ? _T_25942 : 16'h0; // @[Mux.scala 19:72:@20379.4]
  assign _T_25959 = {conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,conflict_9_5,_T_25822}; // @[Mux.scala 19:72:@20394.4]
  assign _T_25961 = _T_2708 ? _T_25959 : 16'h0; // @[Mux.scala 19:72:@20395.4]
  assign _T_25976 = {conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,conflict_9_6,_T_25839}; // @[Mux.scala 19:72:@20410.4]
  assign _T_25978 = _T_2709 ? _T_25976 : 16'h0; // @[Mux.scala 19:72:@20411.4]
  assign _T_25993 = {conflict_9_14,conflict_9_13,conflict_9_12,conflict_9_11,conflict_9_10,conflict_9_9,conflict_9_8,conflict_9_7,_T_25856}; // @[Mux.scala 19:72:@20426.4]
  assign _T_25995 = _T_2710 ? _T_25993 : 16'h0; // @[Mux.scala 19:72:@20427.4]
  assign _T_25996 = _T_25740 | _T_25757; // @[Mux.scala 19:72:@20428.4]
  assign _T_25997 = _T_25996 | _T_25774; // @[Mux.scala 19:72:@20429.4]
  assign _T_25998 = _T_25997 | _T_25791; // @[Mux.scala 19:72:@20430.4]
  assign _T_25999 = _T_25998 | _T_25808; // @[Mux.scala 19:72:@20431.4]
  assign _T_26000 = _T_25999 | _T_25825; // @[Mux.scala 19:72:@20432.4]
  assign _T_26001 = _T_26000 | _T_25842; // @[Mux.scala 19:72:@20433.4]
  assign _T_26002 = _T_26001 | _T_25859; // @[Mux.scala 19:72:@20434.4]
  assign _T_26003 = _T_26002 | _T_25876; // @[Mux.scala 19:72:@20435.4]
  assign _T_26004 = _T_26003 | _T_25893; // @[Mux.scala 19:72:@20436.4]
  assign _T_26005 = _T_26004 | _T_25910; // @[Mux.scala 19:72:@20437.4]
  assign _T_26006 = _T_26005 | _T_25927; // @[Mux.scala 19:72:@20438.4]
  assign _T_26007 = _T_26006 | _T_25944; // @[Mux.scala 19:72:@20439.4]
  assign _T_26008 = _T_26007 | _T_25961; // @[Mux.scala 19:72:@20440.4]
  assign _T_26009 = _T_26008 | _T_25978; // @[Mux.scala 19:72:@20441.4]
  assign _T_26010 = _T_26009 | _T_25995; // @[Mux.scala 19:72:@20442.4]
  assign _T_26588 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0}; // @[Mux.scala 19:72:@20792.4]
  assign _T_26595 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8}; // @[Mux.scala 19:72:@20799.4]
  assign _T_26596 = {conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,_T_26588}; // @[Mux.scala 19:72:@20800.4]
  assign _T_26598 = _T_2695 ? _T_26596 : 16'h0; // @[Mux.scala 19:72:@20801.4]
  assign _T_26605 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1}; // @[Mux.scala 19:72:@20808.4]
  assign _T_26612 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9}; // @[Mux.scala 19:72:@20815.4]
  assign _T_26613 = {conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,_T_26605}; // @[Mux.scala 19:72:@20816.4]
  assign _T_26615 = _T_2696 ? _T_26613 : 16'h0; // @[Mux.scala 19:72:@20817.4]
  assign _T_26622 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2}; // @[Mux.scala 19:72:@20824.4]
  assign _T_26629 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10}; // @[Mux.scala 19:72:@20831.4]
  assign _T_26630 = {conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,_T_26622}; // @[Mux.scala 19:72:@20832.4]
  assign _T_26632 = _T_2697 ? _T_26630 : 16'h0; // @[Mux.scala 19:72:@20833.4]
  assign _T_26639 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3}; // @[Mux.scala 19:72:@20840.4]
  assign _T_26646 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11}; // @[Mux.scala 19:72:@20847.4]
  assign _T_26647 = {conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,_T_26639}; // @[Mux.scala 19:72:@20848.4]
  assign _T_26649 = _T_2698 ? _T_26647 : 16'h0; // @[Mux.scala 19:72:@20849.4]
  assign _T_26656 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4}; // @[Mux.scala 19:72:@20856.4]
  assign _T_26663 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12}; // @[Mux.scala 19:72:@20863.4]
  assign _T_26664 = {conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,conflict_10_12,_T_26656}; // @[Mux.scala 19:72:@20864.4]
  assign _T_26666 = _T_2699 ? _T_26664 : 16'h0; // @[Mux.scala 19:72:@20865.4]
  assign _T_26673 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5}; // @[Mux.scala 19:72:@20872.4]
  assign _T_26680 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13}; // @[Mux.scala 19:72:@20879.4]
  assign _T_26681 = {conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,conflict_10_13,_T_26673}; // @[Mux.scala 19:72:@20880.4]
  assign _T_26683 = _T_2700 ? _T_26681 : 16'h0; // @[Mux.scala 19:72:@20881.4]
  assign _T_26690 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6}; // @[Mux.scala 19:72:@20888.4]
  assign _T_26697 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14}; // @[Mux.scala 19:72:@20895.4]
  assign _T_26698 = {conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,conflict_10_14,_T_26690}; // @[Mux.scala 19:72:@20896.4]
  assign _T_26700 = _T_2701 ? _T_26698 : 16'h0; // @[Mux.scala 19:72:@20897.4]
  assign _T_26707 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7}; // @[Mux.scala 19:72:@20904.4]
  assign _T_26714 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15}; // @[Mux.scala 19:72:@20911.4]
  assign _T_26715 = {conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,conflict_10_15,_T_26707}; // @[Mux.scala 19:72:@20912.4]
  assign _T_26717 = _T_2702 ? _T_26715 : 16'h0; // @[Mux.scala 19:72:@20913.4]
  assign _T_26732 = {conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,conflict_10_0,_T_26595}; // @[Mux.scala 19:72:@20928.4]
  assign _T_26734 = _T_2703 ? _T_26732 : 16'h0; // @[Mux.scala 19:72:@20929.4]
  assign _T_26749 = {conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,conflict_10_1,_T_26612}; // @[Mux.scala 19:72:@20944.4]
  assign _T_26751 = _T_2704 ? _T_26749 : 16'h0; // @[Mux.scala 19:72:@20945.4]
  assign _T_26766 = {conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,conflict_10_2,_T_26629}; // @[Mux.scala 19:72:@20960.4]
  assign _T_26768 = _T_2705 ? _T_26766 : 16'h0; // @[Mux.scala 19:72:@20961.4]
  assign _T_26783 = {conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,conflict_10_3,_T_26646}; // @[Mux.scala 19:72:@20976.4]
  assign _T_26785 = _T_2706 ? _T_26783 : 16'h0; // @[Mux.scala 19:72:@20977.4]
  assign _T_26800 = {conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,conflict_10_4,_T_26663}; // @[Mux.scala 19:72:@20992.4]
  assign _T_26802 = _T_2707 ? _T_26800 : 16'h0; // @[Mux.scala 19:72:@20993.4]
  assign _T_26817 = {conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,conflict_10_5,_T_26680}; // @[Mux.scala 19:72:@21008.4]
  assign _T_26819 = _T_2708 ? _T_26817 : 16'h0; // @[Mux.scala 19:72:@21009.4]
  assign _T_26834 = {conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,conflict_10_6,_T_26697}; // @[Mux.scala 19:72:@21024.4]
  assign _T_26836 = _T_2709 ? _T_26834 : 16'h0; // @[Mux.scala 19:72:@21025.4]
  assign _T_26851 = {conflict_10_14,conflict_10_13,conflict_10_12,conflict_10_11,conflict_10_10,conflict_10_9,conflict_10_8,conflict_10_7,_T_26714}; // @[Mux.scala 19:72:@21040.4]
  assign _T_26853 = _T_2710 ? _T_26851 : 16'h0; // @[Mux.scala 19:72:@21041.4]
  assign _T_26854 = _T_26598 | _T_26615; // @[Mux.scala 19:72:@21042.4]
  assign _T_26855 = _T_26854 | _T_26632; // @[Mux.scala 19:72:@21043.4]
  assign _T_26856 = _T_26855 | _T_26649; // @[Mux.scala 19:72:@21044.4]
  assign _T_26857 = _T_26856 | _T_26666; // @[Mux.scala 19:72:@21045.4]
  assign _T_26858 = _T_26857 | _T_26683; // @[Mux.scala 19:72:@21046.4]
  assign _T_26859 = _T_26858 | _T_26700; // @[Mux.scala 19:72:@21047.4]
  assign _T_26860 = _T_26859 | _T_26717; // @[Mux.scala 19:72:@21048.4]
  assign _T_26861 = _T_26860 | _T_26734; // @[Mux.scala 19:72:@21049.4]
  assign _T_26862 = _T_26861 | _T_26751; // @[Mux.scala 19:72:@21050.4]
  assign _T_26863 = _T_26862 | _T_26768; // @[Mux.scala 19:72:@21051.4]
  assign _T_26864 = _T_26863 | _T_26785; // @[Mux.scala 19:72:@21052.4]
  assign _T_26865 = _T_26864 | _T_26802; // @[Mux.scala 19:72:@21053.4]
  assign _T_26866 = _T_26865 | _T_26819; // @[Mux.scala 19:72:@21054.4]
  assign _T_26867 = _T_26866 | _T_26836; // @[Mux.scala 19:72:@21055.4]
  assign _T_26868 = _T_26867 | _T_26853; // @[Mux.scala 19:72:@21056.4]
  assign _T_27446 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0}; // @[Mux.scala 19:72:@21406.4]
  assign _T_27453 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8}; // @[Mux.scala 19:72:@21413.4]
  assign _T_27454 = {conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,_T_27446}; // @[Mux.scala 19:72:@21414.4]
  assign _T_27456 = _T_2695 ? _T_27454 : 16'h0; // @[Mux.scala 19:72:@21415.4]
  assign _T_27463 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1}; // @[Mux.scala 19:72:@21422.4]
  assign _T_27470 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9}; // @[Mux.scala 19:72:@21429.4]
  assign _T_27471 = {conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,_T_27463}; // @[Mux.scala 19:72:@21430.4]
  assign _T_27473 = _T_2696 ? _T_27471 : 16'h0; // @[Mux.scala 19:72:@21431.4]
  assign _T_27480 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2}; // @[Mux.scala 19:72:@21438.4]
  assign _T_27487 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10}; // @[Mux.scala 19:72:@21445.4]
  assign _T_27488 = {conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,_T_27480}; // @[Mux.scala 19:72:@21446.4]
  assign _T_27490 = _T_2697 ? _T_27488 : 16'h0; // @[Mux.scala 19:72:@21447.4]
  assign _T_27497 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3}; // @[Mux.scala 19:72:@21454.4]
  assign _T_27504 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11}; // @[Mux.scala 19:72:@21461.4]
  assign _T_27505 = {conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,_T_27497}; // @[Mux.scala 19:72:@21462.4]
  assign _T_27507 = _T_2698 ? _T_27505 : 16'h0; // @[Mux.scala 19:72:@21463.4]
  assign _T_27514 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4}; // @[Mux.scala 19:72:@21470.4]
  assign _T_27521 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12}; // @[Mux.scala 19:72:@21477.4]
  assign _T_27522 = {conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,conflict_11_12,_T_27514}; // @[Mux.scala 19:72:@21478.4]
  assign _T_27524 = _T_2699 ? _T_27522 : 16'h0; // @[Mux.scala 19:72:@21479.4]
  assign _T_27531 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5}; // @[Mux.scala 19:72:@21486.4]
  assign _T_27538 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13}; // @[Mux.scala 19:72:@21493.4]
  assign _T_27539 = {conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,conflict_11_13,_T_27531}; // @[Mux.scala 19:72:@21494.4]
  assign _T_27541 = _T_2700 ? _T_27539 : 16'h0; // @[Mux.scala 19:72:@21495.4]
  assign _T_27548 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6}; // @[Mux.scala 19:72:@21502.4]
  assign _T_27555 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14}; // @[Mux.scala 19:72:@21509.4]
  assign _T_27556 = {conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,conflict_11_14,_T_27548}; // @[Mux.scala 19:72:@21510.4]
  assign _T_27558 = _T_2701 ? _T_27556 : 16'h0; // @[Mux.scala 19:72:@21511.4]
  assign _T_27565 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7}; // @[Mux.scala 19:72:@21518.4]
  assign _T_27572 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15}; // @[Mux.scala 19:72:@21525.4]
  assign _T_27573 = {conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,conflict_11_15,_T_27565}; // @[Mux.scala 19:72:@21526.4]
  assign _T_27575 = _T_2702 ? _T_27573 : 16'h0; // @[Mux.scala 19:72:@21527.4]
  assign _T_27590 = {conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,conflict_11_0,_T_27453}; // @[Mux.scala 19:72:@21542.4]
  assign _T_27592 = _T_2703 ? _T_27590 : 16'h0; // @[Mux.scala 19:72:@21543.4]
  assign _T_27607 = {conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,conflict_11_1,_T_27470}; // @[Mux.scala 19:72:@21558.4]
  assign _T_27609 = _T_2704 ? _T_27607 : 16'h0; // @[Mux.scala 19:72:@21559.4]
  assign _T_27624 = {conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,conflict_11_2,_T_27487}; // @[Mux.scala 19:72:@21574.4]
  assign _T_27626 = _T_2705 ? _T_27624 : 16'h0; // @[Mux.scala 19:72:@21575.4]
  assign _T_27641 = {conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,conflict_11_3,_T_27504}; // @[Mux.scala 19:72:@21590.4]
  assign _T_27643 = _T_2706 ? _T_27641 : 16'h0; // @[Mux.scala 19:72:@21591.4]
  assign _T_27658 = {conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,conflict_11_4,_T_27521}; // @[Mux.scala 19:72:@21606.4]
  assign _T_27660 = _T_2707 ? _T_27658 : 16'h0; // @[Mux.scala 19:72:@21607.4]
  assign _T_27675 = {conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,conflict_11_5,_T_27538}; // @[Mux.scala 19:72:@21622.4]
  assign _T_27677 = _T_2708 ? _T_27675 : 16'h0; // @[Mux.scala 19:72:@21623.4]
  assign _T_27692 = {conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,conflict_11_6,_T_27555}; // @[Mux.scala 19:72:@21638.4]
  assign _T_27694 = _T_2709 ? _T_27692 : 16'h0; // @[Mux.scala 19:72:@21639.4]
  assign _T_27709 = {conflict_11_14,conflict_11_13,conflict_11_12,conflict_11_11,conflict_11_10,conflict_11_9,conflict_11_8,conflict_11_7,_T_27572}; // @[Mux.scala 19:72:@21654.4]
  assign _T_27711 = _T_2710 ? _T_27709 : 16'h0; // @[Mux.scala 19:72:@21655.4]
  assign _T_27712 = _T_27456 | _T_27473; // @[Mux.scala 19:72:@21656.4]
  assign _T_27713 = _T_27712 | _T_27490; // @[Mux.scala 19:72:@21657.4]
  assign _T_27714 = _T_27713 | _T_27507; // @[Mux.scala 19:72:@21658.4]
  assign _T_27715 = _T_27714 | _T_27524; // @[Mux.scala 19:72:@21659.4]
  assign _T_27716 = _T_27715 | _T_27541; // @[Mux.scala 19:72:@21660.4]
  assign _T_27717 = _T_27716 | _T_27558; // @[Mux.scala 19:72:@21661.4]
  assign _T_27718 = _T_27717 | _T_27575; // @[Mux.scala 19:72:@21662.4]
  assign _T_27719 = _T_27718 | _T_27592; // @[Mux.scala 19:72:@21663.4]
  assign _T_27720 = _T_27719 | _T_27609; // @[Mux.scala 19:72:@21664.4]
  assign _T_27721 = _T_27720 | _T_27626; // @[Mux.scala 19:72:@21665.4]
  assign _T_27722 = _T_27721 | _T_27643; // @[Mux.scala 19:72:@21666.4]
  assign _T_27723 = _T_27722 | _T_27660; // @[Mux.scala 19:72:@21667.4]
  assign _T_27724 = _T_27723 | _T_27677; // @[Mux.scala 19:72:@21668.4]
  assign _T_27725 = _T_27724 | _T_27694; // @[Mux.scala 19:72:@21669.4]
  assign _T_27726 = _T_27725 | _T_27711; // @[Mux.scala 19:72:@21670.4]
  assign _T_28304 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0}; // @[Mux.scala 19:72:@22020.4]
  assign _T_28311 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8}; // @[Mux.scala 19:72:@22027.4]
  assign _T_28312 = {conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,_T_28304}; // @[Mux.scala 19:72:@22028.4]
  assign _T_28314 = _T_2695 ? _T_28312 : 16'h0; // @[Mux.scala 19:72:@22029.4]
  assign _T_28321 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1}; // @[Mux.scala 19:72:@22036.4]
  assign _T_28328 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9}; // @[Mux.scala 19:72:@22043.4]
  assign _T_28329 = {conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,_T_28321}; // @[Mux.scala 19:72:@22044.4]
  assign _T_28331 = _T_2696 ? _T_28329 : 16'h0; // @[Mux.scala 19:72:@22045.4]
  assign _T_28338 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2}; // @[Mux.scala 19:72:@22052.4]
  assign _T_28345 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10}; // @[Mux.scala 19:72:@22059.4]
  assign _T_28346 = {conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,_T_28338}; // @[Mux.scala 19:72:@22060.4]
  assign _T_28348 = _T_2697 ? _T_28346 : 16'h0; // @[Mux.scala 19:72:@22061.4]
  assign _T_28355 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3}; // @[Mux.scala 19:72:@22068.4]
  assign _T_28362 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11}; // @[Mux.scala 19:72:@22075.4]
  assign _T_28363 = {conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,_T_28355}; // @[Mux.scala 19:72:@22076.4]
  assign _T_28365 = _T_2698 ? _T_28363 : 16'h0; // @[Mux.scala 19:72:@22077.4]
  assign _T_28372 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4}; // @[Mux.scala 19:72:@22084.4]
  assign _T_28379 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12}; // @[Mux.scala 19:72:@22091.4]
  assign _T_28380 = {conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,conflict_12_12,_T_28372}; // @[Mux.scala 19:72:@22092.4]
  assign _T_28382 = _T_2699 ? _T_28380 : 16'h0; // @[Mux.scala 19:72:@22093.4]
  assign _T_28389 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5}; // @[Mux.scala 19:72:@22100.4]
  assign _T_28396 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13}; // @[Mux.scala 19:72:@22107.4]
  assign _T_28397 = {conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,conflict_12_13,_T_28389}; // @[Mux.scala 19:72:@22108.4]
  assign _T_28399 = _T_2700 ? _T_28397 : 16'h0; // @[Mux.scala 19:72:@22109.4]
  assign _T_28406 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6}; // @[Mux.scala 19:72:@22116.4]
  assign _T_28413 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14}; // @[Mux.scala 19:72:@22123.4]
  assign _T_28414 = {conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,conflict_12_14,_T_28406}; // @[Mux.scala 19:72:@22124.4]
  assign _T_28416 = _T_2701 ? _T_28414 : 16'h0; // @[Mux.scala 19:72:@22125.4]
  assign _T_28423 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7}; // @[Mux.scala 19:72:@22132.4]
  assign _T_28430 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15}; // @[Mux.scala 19:72:@22139.4]
  assign _T_28431 = {conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,conflict_12_15,_T_28423}; // @[Mux.scala 19:72:@22140.4]
  assign _T_28433 = _T_2702 ? _T_28431 : 16'h0; // @[Mux.scala 19:72:@22141.4]
  assign _T_28448 = {conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,conflict_12_0,_T_28311}; // @[Mux.scala 19:72:@22156.4]
  assign _T_28450 = _T_2703 ? _T_28448 : 16'h0; // @[Mux.scala 19:72:@22157.4]
  assign _T_28465 = {conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,conflict_12_1,_T_28328}; // @[Mux.scala 19:72:@22172.4]
  assign _T_28467 = _T_2704 ? _T_28465 : 16'h0; // @[Mux.scala 19:72:@22173.4]
  assign _T_28482 = {conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,conflict_12_2,_T_28345}; // @[Mux.scala 19:72:@22188.4]
  assign _T_28484 = _T_2705 ? _T_28482 : 16'h0; // @[Mux.scala 19:72:@22189.4]
  assign _T_28499 = {conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,conflict_12_3,_T_28362}; // @[Mux.scala 19:72:@22204.4]
  assign _T_28501 = _T_2706 ? _T_28499 : 16'h0; // @[Mux.scala 19:72:@22205.4]
  assign _T_28516 = {conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,conflict_12_4,_T_28379}; // @[Mux.scala 19:72:@22220.4]
  assign _T_28518 = _T_2707 ? _T_28516 : 16'h0; // @[Mux.scala 19:72:@22221.4]
  assign _T_28533 = {conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,conflict_12_5,_T_28396}; // @[Mux.scala 19:72:@22236.4]
  assign _T_28535 = _T_2708 ? _T_28533 : 16'h0; // @[Mux.scala 19:72:@22237.4]
  assign _T_28550 = {conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,conflict_12_6,_T_28413}; // @[Mux.scala 19:72:@22252.4]
  assign _T_28552 = _T_2709 ? _T_28550 : 16'h0; // @[Mux.scala 19:72:@22253.4]
  assign _T_28567 = {conflict_12_14,conflict_12_13,conflict_12_12,conflict_12_11,conflict_12_10,conflict_12_9,conflict_12_8,conflict_12_7,_T_28430}; // @[Mux.scala 19:72:@22268.4]
  assign _T_28569 = _T_2710 ? _T_28567 : 16'h0; // @[Mux.scala 19:72:@22269.4]
  assign _T_28570 = _T_28314 | _T_28331; // @[Mux.scala 19:72:@22270.4]
  assign _T_28571 = _T_28570 | _T_28348; // @[Mux.scala 19:72:@22271.4]
  assign _T_28572 = _T_28571 | _T_28365; // @[Mux.scala 19:72:@22272.4]
  assign _T_28573 = _T_28572 | _T_28382; // @[Mux.scala 19:72:@22273.4]
  assign _T_28574 = _T_28573 | _T_28399; // @[Mux.scala 19:72:@22274.4]
  assign _T_28575 = _T_28574 | _T_28416; // @[Mux.scala 19:72:@22275.4]
  assign _T_28576 = _T_28575 | _T_28433; // @[Mux.scala 19:72:@22276.4]
  assign _T_28577 = _T_28576 | _T_28450; // @[Mux.scala 19:72:@22277.4]
  assign _T_28578 = _T_28577 | _T_28467; // @[Mux.scala 19:72:@22278.4]
  assign _T_28579 = _T_28578 | _T_28484; // @[Mux.scala 19:72:@22279.4]
  assign _T_28580 = _T_28579 | _T_28501; // @[Mux.scala 19:72:@22280.4]
  assign _T_28581 = _T_28580 | _T_28518; // @[Mux.scala 19:72:@22281.4]
  assign _T_28582 = _T_28581 | _T_28535; // @[Mux.scala 19:72:@22282.4]
  assign _T_28583 = _T_28582 | _T_28552; // @[Mux.scala 19:72:@22283.4]
  assign _T_28584 = _T_28583 | _T_28569; // @[Mux.scala 19:72:@22284.4]
  assign _T_29162 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0}; // @[Mux.scala 19:72:@22634.4]
  assign _T_29169 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8}; // @[Mux.scala 19:72:@22641.4]
  assign _T_29170 = {conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,_T_29162}; // @[Mux.scala 19:72:@22642.4]
  assign _T_29172 = _T_2695 ? _T_29170 : 16'h0; // @[Mux.scala 19:72:@22643.4]
  assign _T_29179 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1}; // @[Mux.scala 19:72:@22650.4]
  assign _T_29186 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9}; // @[Mux.scala 19:72:@22657.4]
  assign _T_29187 = {conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,_T_29179}; // @[Mux.scala 19:72:@22658.4]
  assign _T_29189 = _T_2696 ? _T_29187 : 16'h0; // @[Mux.scala 19:72:@22659.4]
  assign _T_29196 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2}; // @[Mux.scala 19:72:@22666.4]
  assign _T_29203 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10}; // @[Mux.scala 19:72:@22673.4]
  assign _T_29204 = {conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,_T_29196}; // @[Mux.scala 19:72:@22674.4]
  assign _T_29206 = _T_2697 ? _T_29204 : 16'h0; // @[Mux.scala 19:72:@22675.4]
  assign _T_29213 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3}; // @[Mux.scala 19:72:@22682.4]
  assign _T_29220 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11}; // @[Mux.scala 19:72:@22689.4]
  assign _T_29221 = {conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,_T_29213}; // @[Mux.scala 19:72:@22690.4]
  assign _T_29223 = _T_2698 ? _T_29221 : 16'h0; // @[Mux.scala 19:72:@22691.4]
  assign _T_29230 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4}; // @[Mux.scala 19:72:@22698.4]
  assign _T_29237 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12}; // @[Mux.scala 19:72:@22705.4]
  assign _T_29238 = {conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,conflict_13_12,_T_29230}; // @[Mux.scala 19:72:@22706.4]
  assign _T_29240 = _T_2699 ? _T_29238 : 16'h0; // @[Mux.scala 19:72:@22707.4]
  assign _T_29247 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5}; // @[Mux.scala 19:72:@22714.4]
  assign _T_29254 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13}; // @[Mux.scala 19:72:@22721.4]
  assign _T_29255 = {conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,conflict_13_13,_T_29247}; // @[Mux.scala 19:72:@22722.4]
  assign _T_29257 = _T_2700 ? _T_29255 : 16'h0; // @[Mux.scala 19:72:@22723.4]
  assign _T_29264 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6}; // @[Mux.scala 19:72:@22730.4]
  assign _T_29271 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14}; // @[Mux.scala 19:72:@22737.4]
  assign _T_29272 = {conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,conflict_13_14,_T_29264}; // @[Mux.scala 19:72:@22738.4]
  assign _T_29274 = _T_2701 ? _T_29272 : 16'h0; // @[Mux.scala 19:72:@22739.4]
  assign _T_29281 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7}; // @[Mux.scala 19:72:@22746.4]
  assign _T_29288 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15}; // @[Mux.scala 19:72:@22753.4]
  assign _T_29289 = {conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,conflict_13_15,_T_29281}; // @[Mux.scala 19:72:@22754.4]
  assign _T_29291 = _T_2702 ? _T_29289 : 16'h0; // @[Mux.scala 19:72:@22755.4]
  assign _T_29306 = {conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,conflict_13_0,_T_29169}; // @[Mux.scala 19:72:@22770.4]
  assign _T_29308 = _T_2703 ? _T_29306 : 16'h0; // @[Mux.scala 19:72:@22771.4]
  assign _T_29323 = {conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,conflict_13_1,_T_29186}; // @[Mux.scala 19:72:@22786.4]
  assign _T_29325 = _T_2704 ? _T_29323 : 16'h0; // @[Mux.scala 19:72:@22787.4]
  assign _T_29340 = {conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,conflict_13_2,_T_29203}; // @[Mux.scala 19:72:@22802.4]
  assign _T_29342 = _T_2705 ? _T_29340 : 16'h0; // @[Mux.scala 19:72:@22803.4]
  assign _T_29357 = {conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,conflict_13_3,_T_29220}; // @[Mux.scala 19:72:@22818.4]
  assign _T_29359 = _T_2706 ? _T_29357 : 16'h0; // @[Mux.scala 19:72:@22819.4]
  assign _T_29374 = {conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,conflict_13_4,_T_29237}; // @[Mux.scala 19:72:@22834.4]
  assign _T_29376 = _T_2707 ? _T_29374 : 16'h0; // @[Mux.scala 19:72:@22835.4]
  assign _T_29391 = {conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,conflict_13_5,_T_29254}; // @[Mux.scala 19:72:@22850.4]
  assign _T_29393 = _T_2708 ? _T_29391 : 16'h0; // @[Mux.scala 19:72:@22851.4]
  assign _T_29408 = {conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,conflict_13_6,_T_29271}; // @[Mux.scala 19:72:@22866.4]
  assign _T_29410 = _T_2709 ? _T_29408 : 16'h0; // @[Mux.scala 19:72:@22867.4]
  assign _T_29425 = {conflict_13_14,conflict_13_13,conflict_13_12,conflict_13_11,conflict_13_10,conflict_13_9,conflict_13_8,conflict_13_7,_T_29288}; // @[Mux.scala 19:72:@22882.4]
  assign _T_29427 = _T_2710 ? _T_29425 : 16'h0; // @[Mux.scala 19:72:@22883.4]
  assign _T_29428 = _T_29172 | _T_29189; // @[Mux.scala 19:72:@22884.4]
  assign _T_29429 = _T_29428 | _T_29206; // @[Mux.scala 19:72:@22885.4]
  assign _T_29430 = _T_29429 | _T_29223; // @[Mux.scala 19:72:@22886.4]
  assign _T_29431 = _T_29430 | _T_29240; // @[Mux.scala 19:72:@22887.4]
  assign _T_29432 = _T_29431 | _T_29257; // @[Mux.scala 19:72:@22888.4]
  assign _T_29433 = _T_29432 | _T_29274; // @[Mux.scala 19:72:@22889.4]
  assign _T_29434 = _T_29433 | _T_29291; // @[Mux.scala 19:72:@22890.4]
  assign _T_29435 = _T_29434 | _T_29308; // @[Mux.scala 19:72:@22891.4]
  assign _T_29436 = _T_29435 | _T_29325; // @[Mux.scala 19:72:@22892.4]
  assign _T_29437 = _T_29436 | _T_29342; // @[Mux.scala 19:72:@22893.4]
  assign _T_29438 = _T_29437 | _T_29359; // @[Mux.scala 19:72:@22894.4]
  assign _T_29439 = _T_29438 | _T_29376; // @[Mux.scala 19:72:@22895.4]
  assign _T_29440 = _T_29439 | _T_29393; // @[Mux.scala 19:72:@22896.4]
  assign _T_29441 = _T_29440 | _T_29410; // @[Mux.scala 19:72:@22897.4]
  assign _T_29442 = _T_29441 | _T_29427; // @[Mux.scala 19:72:@22898.4]
  assign _T_30020 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0}; // @[Mux.scala 19:72:@23248.4]
  assign _T_30027 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8}; // @[Mux.scala 19:72:@23255.4]
  assign _T_30028 = {conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,_T_30020}; // @[Mux.scala 19:72:@23256.4]
  assign _T_30030 = _T_2695 ? _T_30028 : 16'h0; // @[Mux.scala 19:72:@23257.4]
  assign _T_30037 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1}; // @[Mux.scala 19:72:@23264.4]
  assign _T_30044 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9}; // @[Mux.scala 19:72:@23271.4]
  assign _T_30045 = {conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,_T_30037}; // @[Mux.scala 19:72:@23272.4]
  assign _T_30047 = _T_2696 ? _T_30045 : 16'h0; // @[Mux.scala 19:72:@23273.4]
  assign _T_30054 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2}; // @[Mux.scala 19:72:@23280.4]
  assign _T_30061 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10}; // @[Mux.scala 19:72:@23287.4]
  assign _T_30062 = {conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,_T_30054}; // @[Mux.scala 19:72:@23288.4]
  assign _T_30064 = _T_2697 ? _T_30062 : 16'h0; // @[Mux.scala 19:72:@23289.4]
  assign _T_30071 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3}; // @[Mux.scala 19:72:@23296.4]
  assign _T_30078 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11}; // @[Mux.scala 19:72:@23303.4]
  assign _T_30079 = {conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,_T_30071}; // @[Mux.scala 19:72:@23304.4]
  assign _T_30081 = _T_2698 ? _T_30079 : 16'h0; // @[Mux.scala 19:72:@23305.4]
  assign _T_30088 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4}; // @[Mux.scala 19:72:@23312.4]
  assign _T_30095 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12}; // @[Mux.scala 19:72:@23319.4]
  assign _T_30096 = {conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,conflict_14_12,_T_30088}; // @[Mux.scala 19:72:@23320.4]
  assign _T_30098 = _T_2699 ? _T_30096 : 16'h0; // @[Mux.scala 19:72:@23321.4]
  assign _T_30105 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5}; // @[Mux.scala 19:72:@23328.4]
  assign _T_30112 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13}; // @[Mux.scala 19:72:@23335.4]
  assign _T_30113 = {conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,conflict_14_13,_T_30105}; // @[Mux.scala 19:72:@23336.4]
  assign _T_30115 = _T_2700 ? _T_30113 : 16'h0; // @[Mux.scala 19:72:@23337.4]
  assign _T_30122 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6}; // @[Mux.scala 19:72:@23344.4]
  assign _T_30129 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14}; // @[Mux.scala 19:72:@23351.4]
  assign _T_30130 = {conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,conflict_14_14,_T_30122}; // @[Mux.scala 19:72:@23352.4]
  assign _T_30132 = _T_2701 ? _T_30130 : 16'h0; // @[Mux.scala 19:72:@23353.4]
  assign _T_30139 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7}; // @[Mux.scala 19:72:@23360.4]
  assign _T_30146 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15}; // @[Mux.scala 19:72:@23367.4]
  assign _T_30147 = {conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,conflict_14_15,_T_30139}; // @[Mux.scala 19:72:@23368.4]
  assign _T_30149 = _T_2702 ? _T_30147 : 16'h0; // @[Mux.scala 19:72:@23369.4]
  assign _T_30164 = {conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,conflict_14_0,_T_30027}; // @[Mux.scala 19:72:@23384.4]
  assign _T_30166 = _T_2703 ? _T_30164 : 16'h0; // @[Mux.scala 19:72:@23385.4]
  assign _T_30181 = {conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,conflict_14_1,_T_30044}; // @[Mux.scala 19:72:@23400.4]
  assign _T_30183 = _T_2704 ? _T_30181 : 16'h0; // @[Mux.scala 19:72:@23401.4]
  assign _T_30198 = {conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,conflict_14_2,_T_30061}; // @[Mux.scala 19:72:@23416.4]
  assign _T_30200 = _T_2705 ? _T_30198 : 16'h0; // @[Mux.scala 19:72:@23417.4]
  assign _T_30215 = {conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,conflict_14_3,_T_30078}; // @[Mux.scala 19:72:@23432.4]
  assign _T_30217 = _T_2706 ? _T_30215 : 16'h0; // @[Mux.scala 19:72:@23433.4]
  assign _T_30232 = {conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,conflict_14_4,_T_30095}; // @[Mux.scala 19:72:@23448.4]
  assign _T_30234 = _T_2707 ? _T_30232 : 16'h0; // @[Mux.scala 19:72:@23449.4]
  assign _T_30249 = {conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,conflict_14_5,_T_30112}; // @[Mux.scala 19:72:@23464.4]
  assign _T_30251 = _T_2708 ? _T_30249 : 16'h0; // @[Mux.scala 19:72:@23465.4]
  assign _T_30266 = {conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,conflict_14_6,_T_30129}; // @[Mux.scala 19:72:@23480.4]
  assign _T_30268 = _T_2709 ? _T_30266 : 16'h0; // @[Mux.scala 19:72:@23481.4]
  assign _T_30283 = {conflict_14_14,conflict_14_13,conflict_14_12,conflict_14_11,conflict_14_10,conflict_14_9,conflict_14_8,conflict_14_7,_T_30146}; // @[Mux.scala 19:72:@23496.4]
  assign _T_30285 = _T_2710 ? _T_30283 : 16'h0; // @[Mux.scala 19:72:@23497.4]
  assign _T_30286 = _T_30030 | _T_30047; // @[Mux.scala 19:72:@23498.4]
  assign _T_30287 = _T_30286 | _T_30064; // @[Mux.scala 19:72:@23499.4]
  assign _T_30288 = _T_30287 | _T_30081; // @[Mux.scala 19:72:@23500.4]
  assign _T_30289 = _T_30288 | _T_30098; // @[Mux.scala 19:72:@23501.4]
  assign _T_30290 = _T_30289 | _T_30115; // @[Mux.scala 19:72:@23502.4]
  assign _T_30291 = _T_30290 | _T_30132; // @[Mux.scala 19:72:@23503.4]
  assign _T_30292 = _T_30291 | _T_30149; // @[Mux.scala 19:72:@23504.4]
  assign _T_30293 = _T_30292 | _T_30166; // @[Mux.scala 19:72:@23505.4]
  assign _T_30294 = _T_30293 | _T_30183; // @[Mux.scala 19:72:@23506.4]
  assign _T_30295 = _T_30294 | _T_30200; // @[Mux.scala 19:72:@23507.4]
  assign _T_30296 = _T_30295 | _T_30217; // @[Mux.scala 19:72:@23508.4]
  assign _T_30297 = _T_30296 | _T_30234; // @[Mux.scala 19:72:@23509.4]
  assign _T_30298 = _T_30297 | _T_30251; // @[Mux.scala 19:72:@23510.4]
  assign _T_30299 = _T_30298 | _T_30268; // @[Mux.scala 19:72:@23511.4]
  assign _T_30300 = _T_30299 | _T_30285; // @[Mux.scala 19:72:@23512.4]
  assign _T_30878 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0}; // @[Mux.scala 19:72:@23862.4]
  assign _T_30885 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8}; // @[Mux.scala 19:72:@23869.4]
  assign _T_30886 = {conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,_T_30878}; // @[Mux.scala 19:72:@23870.4]
  assign _T_30888 = _T_2695 ? _T_30886 : 16'h0; // @[Mux.scala 19:72:@23871.4]
  assign _T_30895 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1}; // @[Mux.scala 19:72:@23878.4]
  assign _T_30902 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9}; // @[Mux.scala 19:72:@23885.4]
  assign _T_30903 = {conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,_T_30895}; // @[Mux.scala 19:72:@23886.4]
  assign _T_30905 = _T_2696 ? _T_30903 : 16'h0; // @[Mux.scala 19:72:@23887.4]
  assign _T_30912 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2}; // @[Mux.scala 19:72:@23894.4]
  assign _T_30919 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10}; // @[Mux.scala 19:72:@23901.4]
  assign _T_30920 = {conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,_T_30912}; // @[Mux.scala 19:72:@23902.4]
  assign _T_30922 = _T_2697 ? _T_30920 : 16'h0; // @[Mux.scala 19:72:@23903.4]
  assign _T_30929 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3}; // @[Mux.scala 19:72:@23910.4]
  assign _T_30936 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11}; // @[Mux.scala 19:72:@23917.4]
  assign _T_30937 = {conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,_T_30929}; // @[Mux.scala 19:72:@23918.4]
  assign _T_30939 = _T_2698 ? _T_30937 : 16'h0; // @[Mux.scala 19:72:@23919.4]
  assign _T_30946 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4}; // @[Mux.scala 19:72:@23926.4]
  assign _T_30953 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12}; // @[Mux.scala 19:72:@23933.4]
  assign _T_30954 = {conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,conflict_15_12,_T_30946}; // @[Mux.scala 19:72:@23934.4]
  assign _T_30956 = _T_2699 ? _T_30954 : 16'h0; // @[Mux.scala 19:72:@23935.4]
  assign _T_30963 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5}; // @[Mux.scala 19:72:@23942.4]
  assign _T_30970 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13}; // @[Mux.scala 19:72:@23949.4]
  assign _T_30971 = {conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,conflict_15_13,_T_30963}; // @[Mux.scala 19:72:@23950.4]
  assign _T_30973 = _T_2700 ? _T_30971 : 16'h0; // @[Mux.scala 19:72:@23951.4]
  assign _T_30980 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6}; // @[Mux.scala 19:72:@23958.4]
  assign _T_30987 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14}; // @[Mux.scala 19:72:@23965.4]
  assign _T_30988 = {conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,conflict_15_14,_T_30980}; // @[Mux.scala 19:72:@23966.4]
  assign _T_30990 = _T_2701 ? _T_30988 : 16'h0; // @[Mux.scala 19:72:@23967.4]
  assign _T_30997 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7}; // @[Mux.scala 19:72:@23974.4]
  assign _T_31004 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15}; // @[Mux.scala 19:72:@23981.4]
  assign _T_31005 = {conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,conflict_15_15,_T_30997}; // @[Mux.scala 19:72:@23982.4]
  assign _T_31007 = _T_2702 ? _T_31005 : 16'h0; // @[Mux.scala 19:72:@23983.4]
  assign _T_31022 = {conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,conflict_15_0,_T_30885}; // @[Mux.scala 19:72:@23998.4]
  assign _T_31024 = _T_2703 ? _T_31022 : 16'h0; // @[Mux.scala 19:72:@23999.4]
  assign _T_31039 = {conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,conflict_15_1,_T_30902}; // @[Mux.scala 19:72:@24014.4]
  assign _T_31041 = _T_2704 ? _T_31039 : 16'h0; // @[Mux.scala 19:72:@24015.4]
  assign _T_31056 = {conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,conflict_15_2,_T_30919}; // @[Mux.scala 19:72:@24030.4]
  assign _T_31058 = _T_2705 ? _T_31056 : 16'h0; // @[Mux.scala 19:72:@24031.4]
  assign _T_31073 = {conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,conflict_15_3,_T_30936}; // @[Mux.scala 19:72:@24046.4]
  assign _T_31075 = _T_2706 ? _T_31073 : 16'h0; // @[Mux.scala 19:72:@24047.4]
  assign _T_31090 = {conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,conflict_15_4,_T_30953}; // @[Mux.scala 19:72:@24062.4]
  assign _T_31092 = _T_2707 ? _T_31090 : 16'h0; // @[Mux.scala 19:72:@24063.4]
  assign _T_31107 = {conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,conflict_15_5,_T_30970}; // @[Mux.scala 19:72:@24078.4]
  assign _T_31109 = _T_2708 ? _T_31107 : 16'h0; // @[Mux.scala 19:72:@24079.4]
  assign _T_31124 = {conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,conflict_15_6,_T_30987}; // @[Mux.scala 19:72:@24094.4]
  assign _T_31126 = _T_2709 ? _T_31124 : 16'h0; // @[Mux.scala 19:72:@24095.4]
  assign _T_31141 = {conflict_15_14,conflict_15_13,conflict_15_12,conflict_15_11,conflict_15_10,conflict_15_9,conflict_15_8,conflict_15_7,_T_31004}; // @[Mux.scala 19:72:@24110.4]
  assign _T_31143 = _T_2710 ? _T_31141 : 16'h0; // @[Mux.scala 19:72:@24111.4]
  assign _T_31144 = _T_30888 | _T_30905; // @[Mux.scala 19:72:@24112.4]
  assign _T_31145 = _T_31144 | _T_30922; // @[Mux.scala 19:72:@24113.4]
  assign _T_31146 = _T_31145 | _T_30939; // @[Mux.scala 19:72:@24114.4]
  assign _T_31147 = _T_31146 | _T_30956; // @[Mux.scala 19:72:@24115.4]
  assign _T_31148 = _T_31147 | _T_30973; // @[Mux.scala 19:72:@24116.4]
  assign _T_31149 = _T_31148 | _T_30990; // @[Mux.scala 19:72:@24117.4]
  assign _T_31150 = _T_31149 | _T_31007; // @[Mux.scala 19:72:@24118.4]
  assign _T_31151 = _T_31150 | _T_31024; // @[Mux.scala 19:72:@24119.4]
  assign _T_31152 = _T_31151 | _T_31041; // @[Mux.scala 19:72:@24120.4]
  assign _T_31153 = _T_31152 | _T_31058; // @[Mux.scala 19:72:@24121.4]
  assign _T_31154 = _T_31153 | _T_31075; // @[Mux.scala 19:72:@24122.4]
  assign _T_31155 = _T_31154 | _T_31092; // @[Mux.scala 19:72:@24123.4]
  assign _T_31156 = _T_31155 | _T_31109; // @[Mux.scala 19:72:@24124.4]
  assign _T_31157 = _T_31156 | _T_31126; // @[Mux.scala 19:72:@24125.4]
  assign _T_31158 = _T_31157 | _T_31143; // @[Mux.scala 19:72:@24126.4]
  assign _T_52332 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0}; // @[Mux.scala 19:72:@24990.4]
  assign _T_52339 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8}; // @[Mux.scala 19:72:@24997.4]
  assign _T_52340 = {storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,_T_52332}; // @[Mux.scala 19:72:@24998.4]
  assign _T_52342 = _T_2695 ? _T_52340 : 16'h0; // @[Mux.scala 19:72:@24999.4]
  assign _T_52349 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1}; // @[Mux.scala 19:72:@25006.4]
  assign _T_52356 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9}; // @[Mux.scala 19:72:@25013.4]
  assign _T_52357 = {storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,_T_52349}; // @[Mux.scala 19:72:@25014.4]
  assign _T_52359 = _T_2696 ? _T_52357 : 16'h0; // @[Mux.scala 19:72:@25015.4]
  assign _T_52366 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2}; // @[Mux.scala 19:72:@25022.4]
  assign _T_52373 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10}; // @[Mux.scala 19:72:@25029.4]
  assign _T_52374 = {storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,_T_52366}; // @[Mux.scala 19:72:@25030.4]
  assign _T_52376 = _T_2697 ? _T_52374 : 16'h0; // @[Mux.scala 19:72:@25031.4]
  assign _T_52383 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3}; // @[Mux.scala 19:72:@25038.4]
  assign _T_52390 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11}; // @[Mux.scala 19:72:@25045.4]
  assign _T_52391 = {storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,_T_52383}; // @[Mux.scala 19:72:@25046.4]
  assign _T_52393 = _T_2698 ? _T_52391 : 16'h0; // @[Mux.scala 19:72:@25047.4]
  assign _T_52400 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4}; // @[Mux.scala 19:72:@25054.4]
  assign _T_52407 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12}; // @[Mux.scala 19:72:@25061.4]
  assign _T_52408 = {storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,_T_52400}; // @[Mux.scala 19:72:@25062.4]
  assign _T_52410 = _T_2699 ? _T_52408 : 16'h0; // @[Mux.scala 19:72:@25063.4]
  assign _T_52417 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5}; // @[Mux.scala 19:72:@25070.4]
  assign _T_52424 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13}; // @[Mux.scala 19:72:@25077.4]
  assign _T_52425 = {storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,_T_52417}; // @[Mux.scala 19:72:@25078.4]
  assign _T_52427 = _T_2700 ? _T_52425 : 16'h0; // @[Mux.scala 19:72:@25079.4]
  assign _T_52434 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6}; // @[Mux.scala 19:72:@25086.4]
  assign _T_52441 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14}; // @[Mux.scala 19:72:@25093.4]
  assign _T_52442 = {storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,storeAddrNotKnownFlags_0_14,_T_52434}; // @[Mux.scala 19:72:@25094.4]
  assign _T_52444 = _T_2701 ? _T_52442 : 16'h0; // @[Mux.scala 19:72:@25095.4]
  assign _T_52451 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7}; // @[Mux.scala 19:72:@25102.4]
  assign _T_52458 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15}; // @[Mux.scala 19:72:@25109.4]
  assign _T_52459 = {storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,storeAddrNotKnownFlags_0_15,_T_52451}; // @[Mux.scala 19:72:@25110.4]
  assign _T_52461 = _T_2702 ? _T_52459 : 16'h0; // @[Mux.scala 19:72:@25111.4]
  assign _T_52476 = {storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,storeAddrNotKnownFlags_0_0,_T_52339}; // @[Mux.scala 19:72:@25126.4]
  assign _T_52478 = _T_2703 ? _T_52476 : 16'h0; // @[Mux.scala 19:72:@25127.4]
  assign _T_52493 = {storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,storeAddrNotKnownFlags_0_1,_T_52356}; // @[Mux.scala 19:72:@25142.4]
  assign _T_52495 = _T_2704 ? _T_52493 : 16'h0; // @[Mux.scala 19:72:@25143.4]
  assign _T_52510 = {storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,storeAddrNotKnownFlags_0_2,_T_52373}; // @[Mux.scala 19:72:@25158.4]
  assign _T_52512 = _T_2705 ? _T_52510 : 16'h0; // @[Mux.scala 19:72:@25159.4]
  assign _T_52527 = {storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,storeAddrNotKnownFlags_0_3,_T_52390}; // @[Mux.scala 19:72:@25174.4]
  assign _T_52529 = _T_2706 ? _T_52527 : 16'h0; // @[Mux.scala 19:72:@25175.4]
  assign _T_52544 = {storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,storeAddrNotKnownFlags_0_4,_T_52407}; // @[Mux.scala 19:72:@25190.4]
  assign _T_52546 = _T_2707 ? _T_52544 : 16'h0; // @[Mux.scala 19:72:@25191.4]
  assign _T_52561 = {storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,storeAddrNotKnownFlags_0_5,_T_52424}; // @[Mux.scala 19:72:@25206.4]
  assign _T_52563 = _T_2708 ? _T_52561 : 16'h0; // @[Mux.scala 19:72:@25207.4]
  assign _T_52578 = {storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,storeAddrNotKnownFlags_0_6,_T_52441}; // @[Mux.scala 19:72:@25222.4]
  assign _T_52580 = _T_2709 ? _T_52578 : 16'h0; // @[Mux.scala 19:72:@25223.4]
  assign _T_52595 = {storeAddrNotKnownFlags_0_14,storeAddrNotKnownFlags_0_13,storeAddrNotKnownFlags_0_12,storeAddrNotKnownFlags_0_11,storeAddrNotKnownFlags_0_10,storeAddrNotKnownFlags_0_9,storeAddrNotKnownFlags_0_8,storeAddrNotKnownFlags_0_7,_T_52458}; // @[Mux.scala 19:72:@25238.4]
  assign _T_52597 = _T_2710 ? _T_52595 : 16'h0; // @[Mux.scala 19:72:@25239.4]
  assign _T_52598 = _T_52342 | _T_52359; // @[Mux.scala 19:72:@25240.4]
  assign _T_52599 = _T_52598 | _T_52376; // @[Mux.scala 19:72:@25241.4]
  assign _T_52600 = _T_52599 | _T_52393; // @[Mux.scala 19:72:@25242.4]
  assign _T_52601 = _T_52600 | _T_52410; // @[Mux.scala 19:72:@25243.4]
  assign _T_52602 = _T_52601 | _T_52427; // @[Mux.scala 19:72:@25244.4]
  assign _T_52603 = _T_52602 | _T_52444; // @[Mux.scala 19:72:@25245.4]
  assign _T_52604 = _T_52603 | _T_52461; // @[Mux.scala 19:72:@25246.4]
  assign _T_52605 = _T_52604 | _T_52478; // @[Mux.scala 19:72:@25247.4]
  assign _T_52606 = _T_52605 | _T_52495; // @[Mux.scala 19:72:@25248.4]
  assign _T_52607 = _T_52606 | _T_52512; // @[Mux.scala 19:72:@25249.4]
  assign _T_52608 = _T_52607 | _T_52529; // @[Mux.scala 19:72:@25250.4]
  assign _T_52609 = _T_52608 | _T_52546; // @[Mux.scala 19:72:@25251.4]
  assign _T_52610 = _T_52609 | _T_52563; // @[Mux.scala 19:72:@25252.4]
  assign _T_52611 = _T_52610 | _T_52580; // @[Mux.scala 19:72:@25253.4]
  assign _T_52612 = _T_52611 | _T_52597; // @[Mux.scala 19:72:@25254.4]
  assign _T_53190 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0}; // @[Mux.scala 19:72:@25604.4]
  assign _T_53197 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8}; // @[Mux.scala 19:72:@25611.4]
  assign _T_53198 = {storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,_T_53190}; // @[Mux.scala 19:72:@25612.4]
  assign _T_53200 = _T_2695 ? _T_53198 : 16'h0; // @[Mux.scala 19:72:@25613.4]
  assign _T_53207 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1}; // @[Mux.scala 19:72:@25620.4]
  assign _T_53214 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9}; // @[Mux.scala 19:72:@25627.4]
  assign _T_53215 = {storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,_T_53207}; // @[Mux.scala 19:72:@25628.4]
  assign _T_53217 = _T_2696 ? _T_53215 : 16'h0; // @[Mux.scala 19:72:@25629.4]
  assign _T_53224 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2}; // @[Mux.scala 19:72:@25636.4]
  assign _T_53231 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10}; // @[Mux.scala 19:72:@25643.4]
  assign _T_53232 = {storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,_T_53224}; // @[Mux.scala 19:72:@25644.4]
  assign _T_53234 = _T_2697 ? _T_53232 : 16'h0; // @[Mux.scala 19:72:@25645.4]
  assign _T_53241 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3}; // @[Mux.scala 19:72:@25652.4]
  assign _T_53248 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11}; // @[Mux.scala 19:72:@25659.4]
  assign _T_53249 = {storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,_T_53241}; // @[Mux.scala 19:72:@25660.4]
  assign _T_53251 = _T_2698 ? _T_53249 : 16'h0; // @[Mux.scala 19:72:@25661.4]
  assign _T_53258 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4}; // @[Mux.scala 19:72:@25668.4]
  assign _T_53265 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12}; // @[Mux.scala 19:72:@25675.4]
  assign _T_53266 = {storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,_T_53258}; // @[Mux.scala 19:72:@25676.4]
  assign _T_53268 = _T_2699 ? _T_53266 : 16'h0; // @[Mux.scala 19:72:@25677.4]
  assign _T_53275 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5}; // @[Mux.scala 19:72:@25684.4]
  assign _T_53282 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13}; // @[Mux.scala 19:72:@25691.4]
  assign _T_53283 = {storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,_T_53275}; // @[Mux.scala 19:72:@25692.4]
  assign _T_53285 = _T_2700 ? _T_53283 : 16'h0; // @[Mux.scala 19:72:@25693.4]
  assign _T_53292 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6}; // @[Mux.scala 19:72:@25700.4]
  assign _T_53299 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14}; // @[Mux.scala 19:72:@25707.4]
  assign _T_53300 = {storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,storeAddrNotKnownFlags_1_14,_T_53292}; // @[Mux.scala 19:72:@25708.4]
  assign _T_53302 = _T_2701 ? _T_53300 : 16'h0; // @[Mux.scala 19:72:@25709.4]
  assign _T_53309 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7}; // @[Mux.scala 19:72:@25716.4]
  assign _T_53316 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15}; // @[Mux.scala 19:72:@25723.4]
  assign _T_53317 = {storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,storeAddrNotKnownFlags_1_15,_T_53309}; // @[Mux.scala 19:72:@25724.4]
  assign _T_53319 = _T_2702 ? _T_53317 : 16'h0; // @[Mux.scala 19:72:@25725.4]
  assign _T_53334 = {storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,storeAddrNotKnownFlags_1_0,_T_53197}; // @[Mux.scala 19:72:@25740.4]
  assign _T_53336 = _T_2703 ? _T_53334 : 16'h0; // @[Mux.scala 19:72:@25741.4]
  assign _T_53351 = {storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,storeAddrNotKnownFlags_1_1,_T_53214}; // @[Mux.scala 19:72:@25756.4]
  assign _T_53353 = _T_2704 ? _T_53351 : 16'h0; // @[Mux.scala 19:72:@25757.4]
  assign _T_53368 = {storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,storeAddrNotKnownFlags_1_2,_T_53231}; // @[Mux.scala 19:72:@25772.4]
  assign _T_53370 = _T_2705 ? _T_53368 : 16'h0; // @[Mux.scala 19:72:@25773.4]
  assign _T_53385 = {storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,storeAddrNotKnownFlags_1_3,_T_53248}; // @[Mux.scala 19:72:@25788.4]
  assign _T_53387 = _T_2706 ? _T_53385 : 16'h0; // @[Mux.scala 19:72:@25789.4]
  assign _T_53402 = {storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,storeAddrNotKnownFlags_1_4,_T_53265}; // @[Mux.scala 19:72:@25804.4]
  assign _T_53404 = _T_2707 ? _T_53402 : 16'h0; // @[Mux.scala 19:72:@25805.4]
  assign _T_53419 = {storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,storeAddrNotKnownFlags_1_5,_T_53282}; // @[Mux.scala 19:72:@25820.4]
  assign _T_53421 = _T_2708 ? _T_53419 : 16'h0; // @[Mux.scala 19:72:@25821.4]
  assign _T_53436 = {storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,storeAddrNotKnownFlags_1_6,_T_53299}; // @[Mux.scala 19:72:@25836.4]
  assign _T_53438 = _T_2709 ? _T_53436 : 16'h0; // @[Mux.scala 19:72:@25837.4]
  assign _T_53453 = {storeAddrNotKnownFlags_1_14,storeAddrNotKnownFlags_1_13,storeAddrNotKnownFlags_1_12,storeAddrNotKnownFlags_1_11,storeAddrNotKnownFlags_1_10,storeAddrNotKnownFlags_1_9,storeAddrNotKnownFlags_1_8,storeAddrNotKnownFlags_1_7,_T_53316}; // @[Mux.scala 19:72:@25852.4]
  assign _T_53455 = _T_2710 ? _T_53453 : 16'h0; // @[Mux.scala 19:72:@25853.4]
  assign _T_53456 = _T_53200 | _T_53217; // @[Mux.scala 19:72:@25854.4]
  assign _T_53457 = _T_53456 | _T_53234; // @[Mux.scala 19:72:@25855.4]
  assign _T_53458 = _T_53457 | _T_53251; // @[Mux.scala 19:72:@25856.4]
  assign _T_53459 = _T_53458 | _T_53268; // @[Mux.scala 19:72:@25857.4]
  assign _T_53460 = _T_53459 | _T_53285; // @[Mux.scala 19:72:@25858.4]
  assign _T_53461 = _T_53460 | _T_53302; // @[Mux.scala 19:72:@25859.4]
  assign _T_53462 = _T_53461 | _T_53319; // @[Mux.scala 19:72:@25860.4]
  assign _T_53463 = _T_53462 | _T_53336; // @[Mux.scala 19:72:@25861.4]
  assign _T_53464 = _T_53463 | _T_53353; // @[Mux.scala 19:72:@25862.4]
  assign _T_53465 = _T_53464 | _T_53370; // @[Mux.scala 19:72:@25863.4]
  assign _T_53466 = _T_53465 | _T_53387; // @[Mux.scala 19:72:@25864.4]
  assign _T_53467 = _T_53466 | _T_53404; // @[Mux.scala 19:72:@25865.4]
  assign _T_53468 = _T_53467 | _T_53421; // @[Mux.scala 19:72:@25866.4]
  assign _T_53469 = _T_53468 | _T_53438; // @[Mux.scala 19:72:@25867.4]
  assign _T_53470 = _T_53469 | _T_53455; // @[Mux.scala 19:72:@25868.4]
  assign _T_54048 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0}; // @[Mux.scala 19:72:@26218.4]
  assign _T_54055 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8}; // @[Mux.scala 19:72:@26225.4]
  assign _T_54056 = {storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,_T_54048}; // @[Mux.scala 19:72:@26226.4]
  assign _T_54058 = _T_2695 ? _T_54056 : 16'h0; // @[Mux.scala 19:72:@26227.4]
  assign _T_54065 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1}; // @[Mux.scala 19:72:@26234.4]
  assign _T_54072 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9}; // @[Mux.scala 19:72:@26241.4]
  assign _T_54073 = {storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,_T_54065}; // @[Mux.scala 19:72:@26242.4]
  assign _T_54075 = _T_2696 ? _T_54073 : 16'h0; // @[Mux.scala 19:72:@26243.4]
  assign _T_54082 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2}; // @[Mux.scala 19:72:@26250.4]
  assign _T_54089 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10}; // @[Mux.scala 19:72:@26257.4]
  assign _T_54090 = {storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,_T_54082}; // @[Mux.scala 19:72:@26258.4]
  assign _T_54092 = _T_2697 ? _T_54090 : 16'h0; // @[Mux.scala 19:72:@26259.4]
  assign _T_54099 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3}; // @[Mux.scala 19:72:@26266.4]
  assign _T_54106 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11}; // @[Mux.scala 19:72:@26273.4]
  assign _T_54107 = {storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,_T_54099}; // @[Mux.scala 19:72:@26274.4]
  assign _T_54109 = _T_2698 ? _T_54107 : 16'h0; // @[Mux.scala 19:72:@26275.4]
  assign _T_54116 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4}; // @[Mux.scala 19:72:@26282.4]
  assign _T_54123 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12}; // @[Mux.scala 19:72:@26289.4]
  assign _T_54124 = {storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,_T_54116}; // @[Mux.scala 19:72:@26290.4]
  assign _T_54126 = _T_2699 ? _T_54124 : 16'h0; // @[Mux.scala 19:72:@26291.4]
  assign _T_54133 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5}; // @[Mux.scala 19:72:@26298.4]
  assign _T_54140 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13}; // @[Mux.scala 19:72:@26305.4]
  assign _T_54141 = {storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,_T_54133}; // @[Mux.scala 19:72:@26306.4]
  assign _T_54143 = _T_2700 ? _T_54141 : 16'h0; // @[Mux.scala 19:72:@26307.4]
  assign _T_54150 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6}; // @[Mux.scala 19:72:@26314.4]
  assign _T_54157 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14}; // @[Mux.scala 19:72:@26321.4]
  assign _T_54158 = {storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,storeAddrNotKnownFlags_2_14,_T_54150}; // @[Mux.scala 19:72:@26322.4]
  assign _T_54160 = _T_2701 ? _T_54158 : 16'h0; // @[Mux.scala 19:72:@26323.4]
  assign _T_54167 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7}; // @[Mux.scala 19:72:@26330.4]
  assign _T_54174 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15}; // @[Mux.scala 19:72:@26337.4]
  assign _T_54175 = {storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,storeAddrNotKnownFlags_2_15,_T_54167}; // @[Mux.scala 19:72:@26338.4]
  assign _T_54177 = _T_2702 ? _T_54175 : 16'h0; // @[Mux.scala 19:72:@26339.4]
  assign _T_54192 = {storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,storeAddrNotKnownFlags_2_0,_T_54055}; // @[Mux.scala 19:72:@26354.4]
  assign _T_54194 = _T_2703 ? _T_54192 : 16'h0; // @[Mux.scala 19:72:@26355.4]
  assign _T_54209 = {storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,storeAddrNotKnownFlags_2_1,_T_54072}; // @[Mux.scala 19:72:@26370.4]
  assign _T_54211 = _T_2704 ? _T_54209 : 16'h0; // @[Mux.scala 19:72:@26371.4]
  assign _T_54226 = {storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,storeAddrNotKnownFlags_2_2,_T_54089}; // @[Mux.scala 19:72:@26386.4]
  assign _T_54228 = _T_2705 ? _T_54226 : 16'h0; // @[Mux.scala 19:72:@26387.4]
  assign _T_54243 = {storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,storeAddrNotKnownFlags_2_3,_T_54106}; // @[Mux.scala 19:72:@26402.4]
  assign _T_54245 = _T_2706 ? _T_54243 : 16'h0; // @[Mux.scala 19:72:@26403.4]
  assign _T_54260 = {storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,storeAddrNotKnownFlags_2_4,_T_54123}; // @[Mux.scala 19:72:@26418.4]
  assign _T_54262 = _T_2707 ? _T_54260 : 16'h0; // @[Mux.scala 19:72:@26419.4]
  assign _T_54277 = {storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,storeAddrNotKnownFlags_2_5,_T_54140}; // @[Mux.scala 19:72:@26434.4]
  assign _T_54279 = _T_2708 ? _T_54277 : 16'h0; // @[Mux.scala 19:72:@26435.4]
  assign _T_54294 = {storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,storeAddrNotKnownFlags_2_6,_T_54157}; // @[Mux.scala 19:72:@26450.4]
  assign _T_54296 = _T_2709 ? _T_54294 : 16'h0; // @[Mux.scala 19:72:@26451.4]
  assign _T_54311 = {storeAddrNotKnownFlags_2_14,storeAddrNotKnownFlags_2_13,storeAddrNotKnownFlags_2_12,storeAddrNotKnownFlags_2_11,storeAddrNotKnownFlags_2_10,storeAddrNotKnownFlags_2_9,storeAddrNotKnownFlags_2_8,storeAddrNotKnownFlags_2_7,_T_54174}; // @[Mux.scala 19:72:@26466.4]
  assign _T_54313 = _T_2710 ? _T_54311 : 16'h0; // @[Mux.scala 19:72:@26467.4]
  assign _T_54314 = _T_54058 | _T_54075; // @[Mux.scala 19:72:@26468.4]
  assign _T_54315 = _T_54314 | _T_54092; // @[Mux.scala 19:72:@26469.4]
  assign _T_54316 = _T_54315 | _T_54109; // @[Mux.scala 19:72:@26470.4]
  assign _T_54317 = _T_54316 | _T_54126; // @[Mux.scala 19:72:@26471.4]
  assign _T_54318 = _T_54317 | _T_54143; // @[Mux.scala 19:72:@26472.4]
  assign _T_54319 = _T_54318 | _T_54160; // @[Mux.scala 19:72:@26473.4]
  assign _T_54320 = _T_54319 | _T_54177; // @[Mux.scala 19:72:@26474.4]
  assign _T_54321 = _T_54320 | _T_54194; // @[Mux.scala 19:72:@26475.4]
  assign _T_54322 = _T_54321 | _T_54211; // @[Mux.scala 19:72:@26476.4]
  assign _T_54323 = _T_54322 | _T_54228; // @[Mux.scala 19:72:@26477.4]
  assign _T_54324 = _T_54323 | _T_54245; // @[Mux.scala 19:72:@26478.4]
  assign _T_54325 = _T_54324 | _T_54262; // @[Mux.scala 19:72:@26479.4]
  assign _T_54326 = _T_54325 | _T_54279; // @[Mux.scala 19:72:@26480.4]
  assign _T_54327 = _T_54326 | _T_54296; // @[Mux.scala 19:72:@26481.4]
  assign _T_54328 = _T_54327 | _T_54313; // @[Mux.scala 19:72:@26482.4]
  assign _T_54906 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0}; // @[Mux.scala 19:72:@26832.4]
  assign _T_54913 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8}; // @[Mux.scala 19:72:@26839.4]
  assign _T_54914 = {storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,_T_54906}; // @[Mux.scala 19:72:@26840.4]
  assign _T_54916 = _T_2695 ? _T_54914 : 16'h0; // @[Mux.scala 19:72:@26841.4]
  assign _T_54923 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1}; // @[Mux.scala 19:72:@26848.4]
  assign _T_54930 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9}; // @[Mux.scala 19:72:@26855.4]
  assign _T_54931 = {storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,_T_54923}; // @[Mux.scala 19:72:@26856.4]
  assign _T_54933 = _T_2696 ? _T_54931 : 16'h0; // @[Mux.scala 19:72:@26857.4]
  assign _T_54940 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2}; // @[Mux.scala 19:72:@26864.4]
  assign _T_54947 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10}; // @[Mux.scala 19:72:@26871.4]
  assign _T_54948 = {storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,_T_54940}; // @[Mux.scala 19:72:@26872.4]
  assign _T_54950 = _T_2697 ? _T_54948 : 16'h0; // @[Mux.scala 19:72:@26873.4]
  assign _T_54957 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3}; // @[Mux.scala 19:72:@26880.4]
  assign _T_54964 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11}; // @[Mux.scala 19:72:@26887.4]
  assign _T_54965 = {storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,_T_54957}; // @[Mux.scala 19:72:@26888.4]
  assign _T_54967 = _T_2698 ? _T_54965 : 16'h0; // @[Mux.scala 19:72:@26889.4]
  assign _T_54974 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4}; // @[Mux.scala 19:72:@26896.4]
  assign _T_54981 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12}; // @[Mux.scala 19:72:@26903.4]
  assign _T_54982 = {storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,_T_54974}; // @[Mux.scala 19:72:@26904.4]
  assign _T_54984 = _T_2699 ? _T_54982 : 16'h0; // @[Mux.scala 19:72:@26905.4]
  assign _T_54991 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5}; // @[Mux.scala 19:72:@26912.4]
  assign _T_54998 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13}; // @[Mux.scala 19:72:@26919.4]
  assign _T_54999 = {storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,_T_54991}; // @[Mux.scala 19:72:@26920.4]
  assign _T_55001 = _T_2700 ? _T_54999 : 16'h0; // @[Mux.scala 19:72:@26921.4]
  assign _T_55008 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6}; // @[Mux.scala 19:72:@26928.4]
  assign _T_55015 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14}; // @[Mux.scala 19:72:@26935.4]
  assign _T_55016 = {storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,storeAddrNotKnownFlags_3_14,_T_55008}; // @[Mux.scala 19:72:@26936.4]
  assign _T_55018 = _T_2701 ? _T_55016 : 16'h0; // @[Mux.scala 19:72:@26937.4]
  assign _T_55025 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7}; // @[Mux.scala 19:72:@26944.4]
  assign _T_55032 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15}; // @[Mux.scala 19:72:@26951.4]
  assign _T_55033 = {storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,storeAddrNotKnownFlags_3_15,_T_55025}; // @[Mux.scala 19:72:@26952.4]
  assign _T_55035 = _T_2702 ? _T_55033 : 16'h0; // @[Mux.scala 19:72:@26953.4]
  assign _T_55050 = {storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,storeAddrNotKnownFlags_3_0,_T_54913}; // @[Mux.scala 19:72:@26968.4]
  assign _T_55052 = _T_2703 ? _T_55050 : 16'h0; // @[Mux.scala 19:72:@26969.4]
  assign _T_55067 = {storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,storeAddrNotKnownFlags_3_1,_T_54930}; // @[Mux.scala 19:72:@26984.4]
  assign _T_55069 = _T_2704 ? _T_55067 : 16'h0; // @[Mux.scala 19:72:@26985.4]
  assign _T_55084 = {storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,storeAddrNotKnownFlags_3_2,_T_54947}; // @[Mux.scala 19:72:@27000.4]
  assign _T_55086 = _T_2705 ? _T_55084 : 16'h0; // @[Mux.scala 19:72:@27001.4]
  assign _T_55101 = {storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,storeAddrNotKnownFlags_3_3,_T_54964}; // @[Mux.scala 19:72:@27016.4]
  assign _T_55103 = _T_2706 ? _T_55101 : 16'h0; // @[Mux.scala 19:72:@27017.4]
  assign _T_55118 = {storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,storeAddrNotKnownFlags_3_4,_T_54981}; // @[Mux.scala 19:72:@27032.4]
  assign _T_55120 = _T_2707 ? _T_55118 : 16'h0; // @[Mux.scala 19:72:@27033.4]
  assign _T_55135 = {storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,storeAddrNotKnownFlags_3_5,_T_54998}; // @[Mux.scala 19:72:@27048.4]
  assign _T_55137 = _T_2708 ? _T_55135 : 16'h0; // @[Mux.scala 19:72:@27049.4]
  assign _T_55152 = {storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,storeAddrNotKnownFlags_3_6,_T_55015}; // @[Mux.scala 19:72:@27064.4]
  assign _T_55154 = _T_2709 ? _T_55152 : 16'h0; // @[Mux.scala 19:72:@27065.4]
  assign _T_55169 = {storeAddrNotKnownFlags_3_14,storeAddrNotKnownFlags_3_13,storeAddrNotKnownFlags_3_12,storeAddrNotKnownFlags_3_11,storeAddrNotKnownFlags_3_10,storeAddrNotKnownFlags_3_9,storeAddrNotKnownFlags_3_8,storeAddrNotKnownFlags_3_7,_T_55032}; // @[Mux.scala 19:72:@27080.4]
  assign _T_55171 = _T_2710 ? _T_55169 : 16'h0; // @[Mux.scala 19:72:@27081.4]
  assign _T_55172 = _T_54916 | _T_54933; // @[Mux.scala 19:72:@27082.4]
  assign _T_55173 = _T_55172 | _T_54950; // @[Mux.scala 19:72:@27083.4]
  assign _T_55174 = _T_55173 | _T_54967; // @[Mux.scala 19:72:@27084.4]
  assign _T_55175 = _T_55174 | _T_54984; // @[Mux.scala 19:72:@27085.4]
  assign _T_55176 = _T_55175 | _T_55001; // @[Mux.scala 19:72:@27086.4]
  assign _T_55177 = _T_55176 | _T_55018; // @[Mux.scala 19:72:@27087.4]
  assign _T_55178 = _T_55177 | _T_55035; // @[Mux.scala 19:72:@27088.4]
  assign _T_55179 = _T_55178 | _T_55052; // @[Mux.scala 19:72:@27089.4]
  assign _T_55180 = _T_55179 | _T_55069; // @[Mux.scala 19:72:@27090.4]
  assign _T_55181 = _T_55180 | _T_55086; // @[Mux.scala 19:72:@27091.4]
  assign _T_55182 = _T_55181 | _T_55103; // @[Mux.scala 19:72:@27092.4]
  assign _T_55183 = _T_55182 | _T_55120; // @[Mux.scala 19:72:@27093.4]
  assign _T_55184 = _T_55183 | _T_55137; // @[Mux.scala 19:72:@27094.4]
  assign _T_55185 = _T_55184 | _T_55154; // @[Mux.scala 19:72:@27095.4]
  assign _T_55186 = _T_55185 | _T_55171; // @[Mux.scala 19:72:@27096.4]
  assign _T_55764 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0}; // @[Mux.scala 19:72:@27446.4]
  assign _T_55771 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8}; // @[Mux.scala 19:72:@27453.4]
  assign _T_55772 = {storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,_T_55764}; // @[Mux.scala 19:72:@27454.4]
  assign _T_55774 = _T_2695 ? _T_55772 : 16'h0; // @[Mux.scala 19:72:@27455.4]
  assign _T_55781 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1}; // @[Mux.scala 19:72:@27462.4]
  assign _T_55788 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9}; // @[Mux.scala 19:72:@27469.4]
  assign _T_55789 = {storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,_T_55781}; // @[Mux.scala 19:72:@27470.4]
  assign _T_55791 = _T_2696 ? _T_55789 : 16'h0; // @[Mux.scala 19:72:@27471.4]
  assign _T_55798 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2}; // @[Mux.scala 19:72:@27478.4]
  assign _T_55805 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10}; // @[Mux.scala 19:72:@27485.4]
  assign _T_55806 = {storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,_T_55798}; // @[Mux.scala 19:72:@27486.4]
  assign _T_55808 = _T_2697 ? _T_55806 : 16'h0; // @[Mux.scala 19:72:@27487.4]
  assign _T_55815 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3}; // @[Mux.scala 19:72:@27494.4]
  assign _T_55822 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11}; // @[Mux.scala 19:72:@27501.4]
  assign _T_55823 = {storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,_T_55815}; // @[Mux.scala 19:72:@27502.4]
  assign _T_55825 = _T_2698 ? _T_55823 : 16'h0; // @[Mux.scala 19:72:@27503.4]
  assign _T_55832 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4}; // @[Mux.scala 19:72:@27510.4]
  assign _T_55839 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12}; // @[Mux.scala 19:72:@27517.4]
  assign _T_55840 = {storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,_T_55832}; // @[Mux.scala 19:72:@27518.4]
  assign _T_55842 = _T_2699 ? _T_55840 : 16'h0; // @[Mux.scala 19:72:@27519.4]
  assign _T_55849 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5}; // @[Mux.scala 19:72:@27526.4]
  assign _T_55856 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13}; // @[Mux.scala 19:72:@27533.4]
  assign _T_55857 = {storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,_T_55849}; // @[Mux.scala 19:72:@27534.4]
  assign _T_55859 = _T_2700 ? _T_55857 : 16'h0; // @[Mux.scala 19:72:@27535.4]
  assign _T_55866 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6}; // @[Mux.scala 19:72:@27542.4]
  assign _T_55873 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14}; // @[Mux.scala 19:72:@27549.4]
  assign _T_55874 = {storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,storeAddrNotKnownFlags_4_14,_T_55866}; // @[Mux.scala 19:72:@27550.4]
  assign _T_55876 = _T_2701 ? _T_55874 : 16'h0; // @[Mux.scala 19:72:@27551.4]
  assign _T_55883 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7}; // @[Mux.scala 19:72:@27558.4]
  assign _T_55890 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15}; // @[Mux.scala 19:72:@27565.4]
  assign _T_55891 = {storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,storeAddrNotKnownFlags_4_15,_T_55883}; // @[Mux.scala 19:72:@27566.4]
  assign _T_55893 = _T_2702 ? _T_55891 : 16'h0; // @[Mux.scala 19:72:@27567.4]
  assign _T_55908 = {storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,storeAddrNotKnownFlags_4_0,_T_55771}; // @[Mux.scala 19:72:@27582.4]
  assign _T_55910 = _T_2703 ? _T_55908 : 16'h0; // @[Mux.scala 19:72:@27583.4]
  assign _T_55925 = {storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,storeAddrNotKnownFlags_4_1,_T_55788}; // @[Mux.scala 19:72:@27598.4]
  assign _T_55927 = _T_2704 ? _T_55925 : 16'h0; // @[Mux.scala 19:72:@27599.4]
  assign _T_55942 = {storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,storeAddrNotKnownFlags_4_2,_T_55805}; // @[Mux.scala 19:72:@27614.4]
  assign _T_55944 = _T_2705 ? _T_55942 : 16'h0; // @[Mux.scala 19:72:@27615.4]
  assign _T_55959 = {storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,storeAddrNotKnownFlags_4_3,_T_55822}; // @[Mux.scala 19:72:@27630.4]
  assign _T_55961 = _T_2706 ? _T_55959 : 16'h0; // @[Mux.scala 19:72:@27631.4]
  assign _T_55976 = {storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,storeAddrNotKnownFlags_4_4,_T_55839}; // @[Mux.scala 19:72:@27646.4]
  assign _T_55978 = _T_2707 ? _T_55976 : 16'h0; // @[Mux.scala 19:72:@27647.4]
  assign _T_55993 = {storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,storeAddrNotKnownFlags_4_5,_T_55856}; // @[Mux.scala 19:72:@27662.4]
  assign _T_55995 = _T_2708 ? _T_55993 : 16'h0; // @[Mux.scala 19:72:@27663.4]
  assign _T_56010 = {storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,storeAddrNotKnownFlags_4_6,_T_55873}; // @[Mux.scala 19:72:@27678.4]
  assign _T_56012 = _T_2709 ? _T_56010 : 16'h0; // @[Mux.scala 19:72:@27679.4]
  assign _T_56027 = {storeAddrNotKnownFlags_4_14,storeAddrNotKnownFlags_4_13,storeAddrNotKnownFlags_4_12,storeAddrNotKnownFlags_4_11,storeAddrNotKnownFlags_4_10,storeAddrNotKnownFlags_4_9,storeAddrNotKnownFlags_4_8,storeAddrNotKnownFlags_4_7,_T_55890}; // @[Mux.scala 19:72:@27694.4]
  assign _T_56029 = _T_2710 ? _T_56027 : 16'h0; // @[Mux.scala 19:72:@27695.4]
  assign _T_56030 = _T_55774 | _T_55791; // @[Mux.scala 19:72:@27696.4]
  assign _T_56031 = _T_56030 | _T_55808; // @[Mux.scala 19:72:@27697.4]
  assign _T_56032 = _T_56031 | _T_55825; // @[Mux.scala 19:72:@27698.4]
  assign _T_56033 = _T_56032 | _T_55842; // @[Mux.scala 19:72:@27699.4]
  assign _T_56034 = _T_56033 | _T_55859; // @[Mux.scala 19:72:@27700.4]
  assign _T_56035 = _T_56034 | _T_55876; // @[Mux.scala 19:72:@27701.4]
  assign _T_56036 = _T_56035 | _T_55893; // @[Mux.scala 19:72:@27702.4]
  assign _T_56037 = _T_56036 | _T_55910; // @[Mux.scala 19:72:@27703.4]
  assign _T_56038 = _T_56037 | _T_55927; // @[Mux.scala 19:72:@27704.4]
  assign _T_56039 = _T_56038 | _T_55944; // @[Mux.scala 19:72:@27705.4]
  assign _T_56040 = _T_56039 | _T_55961; // @[Mux.scala 19:72:@27706.4]
  assign _T_56041 = _T_56040 | _T_55978; // @[Mux.scala 19:72:@27707.4]
  assign _T_56042 = _T_56041 | _T_55995; // @[Mux.scala 19:72:@27708.4]
  assign _T_56043 = _T_56042 | _T_56012; // @[Mux.scala 19:72:@27709.4]
  assign _T_56044 = _T_56043 | _T_56029; // @[Mux.scala 19:72:@27710.4]
  assign _T_56622 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0}; // @[Mux.scala 19:72:@28060.4]
  assign _T_56629 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8}; // @[Mux.scala 19:72:@28067.4]
  assign _T_56630 = {storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,_T_56622}; // @[Mux.scala 19:72:@28068.4]
  assign _T_56632 = _T_2695 ? _T_56630 : 16'h0; // @[Mux.scala 19:72:@28069.4]
  assign _T_56639 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1}; // @[Mux.scala 19:72:@28076.4]
  assign _T_56646 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9}; // @[Mux.scala 19:72:@28083.4]
  assign _T_56647 = {storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,_T_56639}; // @[Mux.scala 19:72:@28084.4]
  assign _T_56649 = _T_2696 ? _T_56647 : 16'h0; // @[Mux.scala 19:72:@28085.4]
  assign _T_56656 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2}; // @[Mux.scala 19:72:@28092.4]
  assign _T_56663 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10}; // @[Mux.scala 19:72:@28099.4]
  assign _T_56664 = {storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,_T_56656}; // @[Mux.scala 19:72:@28100.4]
  assign _T_56666 = _T_2697 ? _T_56664 : 16'h0; // @[Mux.scala 19:72:@28101.4]
  assign _T_56673 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3}; // @[Mux.scala 19:72:@28108.4]
  assign _T_56680 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11}; // @[Mux.scala 19:72:@28115.4]
  assign _T_56681 = {storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,_T_56673}; // @[Mux.scala 19:72:@28116.4]
  assign _T_56683 = _T_2698 ? _T_56681 : 16'h0; // @[Mux.scala 19:72:@28117.4]
  assign _T_56690 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4}; // @[Mux.scala 19:72:@28124.4]
  assign _T_56697 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12}; // @[Mux.scala 19:72:@28131.4]
  assign _T_56698 = {storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,_T_56690}; // @[Mux.scala 19:72:@28132.4]
  assign _T_56700 = _T_2699 ? _T_56698 : 16'h0; // @[Mux.scala 19:72:@28133.4]
  assign _T_56707 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5}; // @[Mux.scala 19:72:@28140.4]
  assign _T_56714 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13}; // @[Mux.scala 19:72:@28147.4]
  assign _T_56715 = {storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,_T_56707}; // @[Mux.scala 19:72:@28148.4]
  assign _T_56717 = _T_2700 ? _T_56715 : 16'h0; // @[Mux.scala 19:72:@28149.4]
  assign _T_56724 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6}; // @[Mux.scala 19:72:@28156.4]
  assign _T_56731 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14}; // @[Mux.scala 19:72:@28163.4]
  assign _T_56732 = {storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,storeAddrNotKnownFlags_5_14,_T_56724}; // @[Mux.scala 19:72:@28164.4]
  assign _T_56734 = _T_2701 ? _T_56732 : 16'h0; // @[Mux.scala 19:72:@28165.4]
  assign _T_56741 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7}; // @[Mux.scala 19:72:@28172.4]
  assign _T_56748 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15}; // @[Mux.scala 19:72:@28179.4]
  assign _T_56749 = {storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,storeAddrNotKnownFlags_5_15,_T_56741}; // @[Mux.scala 19:72:@28180.4]
  assign _T_56751 = _T_2702 ? _T_56749 : 16'h0; // @[Mux.scala 19:72:@28181.4]
  assign _T_56766 = {storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,storeAddrNotKnownFlags_5_0,_T_56629}; // @[Mux.scala 19:72:@28196.4]
  assign _T_56768 = _T_2703 ? _T_56766 : 16'h0; // @[Mux.scala 19:72:@28197.4]
  assign _T_56783 = {storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,storeAddrNotKnownFlags_5_1,_T_56646}; // @[Mux.scala 19:72:@28212.4]
  assign _T_56785 = _T_2704 ? _T_56783 : 16'h0; // @[Mux.scala 19:72:@28213.4]
  assign _T_56800 = {storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,storeAddrNotKnownFlags_5_2,_T_56663}; // @[Mux.scala 19:72:@28228.4]
  assign _T_56802 = _T_2705 ? _T_56800 : 16'h0; // @[Mux.scala 19:72:@28229.4]
  assign _T_56817 = {storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,storeAddrNotKnownFlags_5_3,_T_56680}; // @[Mux.scala 19:72:@28244.4]
  assign _T_56819 = _T_2706 ? _T_56817 : 16'h0; // @[Mux.scala 19:72:@28245.4]
  assign _T_56834 = {storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,storeAddrNotKnownFlags_5_4,_T_56697}; // @[Mux.scala 19:72:@28260.4]
  assign _T_56836 = _T_2707 ? _T_56834 : 16'h0; // @[Mux.scala 19:72:@28261.4]
  assign _T_56851 = {storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,storeAddrNotKnownFlags_5_5,_T_56714}; // @[Mux.scala 19:72:@28276.4]
  assign _T_56853 = _T_2708 ? _T_56851 : 16'h0; // @[Mux.scala 19:72:@28277.4]
  assign _T_56868 = {storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,storeAddrNotKnownFlags_5_6,_T_56731}; // @[Mux.scala 19:72:@28292.4]
  assign _T_56870 = _T_2709 ? _T_56868 : 16'h0; // @[Mux.scala 19:72:@28293.4]
  assign _T_56885 = {storeAddrNotKnownFlags_5_14,storeAddrNotKnownFlags_5_13,storeAddrNotKnownFlags_5_12,storeAddrNotKnownFlags_5_11,storeAddrNotKnownFlags_5_10,storeAddrNotKnownFlags_5_9,storeAddrNotKnownFlags_5_8,storeAddrNotKnownFlags_5_7,_T_56748}; // @[Mux.scala 19:72:@28308.4]
  assign _T_56887 = _T_2710 ? _T_56885 : 16'h0; // @[Mux.scala 19:72:@28309.4]
  assign _T_56888 = _T_56632 | _T_56649; // @[Mux.scala 19:72:@28310.4]
  assign _T_56889 = _T_56888 | _T_56666; // @[Mux.scala 19:72:@28311.4]
  assign _T_56890 = _T_56889 | _T_56683; // @[Mux.scala 19:72:@28312.4]
  assign _T_56891 = _T_56890 | _T_56700; // @[Mux.scala 19:72:@28313.4]
  assign _T_56892 = _T_56891 | _T_56717; // @[Mux.scala 19:72:@28314.4]
  assign _T_56893 = _T_56892 | _T_56734; // @[Mux.scala 19:72:@28315.4]
  assign _T_56894 = _T_56893 | _T_56751; // @[Mux.scala 19:72:@28316.4]
  assign _T_56895 = _T_56894 | _T_56768; // @[Mux.scala 19:72:@28317.4]
  assign _T_56896 = _T_56895 | _T_56785; // @[Mux.scala 19:72:@28318.4]
  assign _T_56897 = _T_56896 | _T_56802; // @[Mux.scala 19:72:@28319.4]
  assign _T_56898 = _T_56897 | _T_56819; // @[Mux.scala 19:72:@28320.4]
  assign _T_56899 = _T_56898 | _T_56836; // @[Mux.scala 19:72:@28321.4]
  assign _T_56900 = _T_56899 | _T_56853; // @[Mux.scala 19:72:@28322.4]
  assign _T_56901 = _T_56900 | _T_56870; // @[Mux.scala 19:72:@28323.4]
  assign _T_56902 = _T_56901 | _T_56887; // @[Mux.scala 19:72:@28324.4]
  assign _T_57480 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0}; // @[Mux.scala 19:72:@28674.4]
  assign _T_57487 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8}; // @[Mux.scala 19:72:@28681.4]
  assign _T_57488 = {storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,_T_57480}; // @[Mux.scala 19:72:@28682.4]
  assign _T_57490 = _T_2695 ? _T_57488 : 16'h0; // @[Mux.scala 19:72:@28683.4]
  assign _T_57497 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1}; // @[Mux.scala 19:72:@28690.4]
  assign _T_57504 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9}; // @[Mux.scala 19:72:@28697.4]
  assign _T_57505 = {storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,_T_57497}; // @[Mux.scala 19:72:@28698.4]
  assign _T_57507 = _T_2696 ? _T_57505 : 16'h0; // @[Mux.scala 19:72:@28699.4]
  assign _T_57514 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2}; // @[Mux.scala 19:72:@28706.4]
  assign _T_57521 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10}; // @[Mux.scala 19:72:@28713.4]
  assign _T_57522 = {storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,_T_57514}; // @[Mux.scala 19:72:@28714.4]
  assign _T_57524 = _T_2697 ? _T_57522 : 16'h0; // @[Mux.scala 19:72:@28715.4]
  assign _T_57531 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3}; // @[Mux.scala 19:72:@28722.4]
  assign _T_57538 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11}; // @[Mux.scala 19:72:@28729.4]
  assign _T_57539 = {storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,_T_57531}; // @[Mux.scala 19:72:@28730.4]
  assign _T_57541 = _T_2698 ? _T_57539 : 16'h0; // @[Mux.scala 19:72:@28731.4]
  assign _T_57548 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4}; // @[Mux.scala 19:72:@28738.4]
  assign _T_57555 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12}; // @[Mux.scala 19:72:@28745.4]
  assign _T_57556 = {storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,_T_57548}; // @[Mux.scala 19:72:@28746.4]
  assign _T_57558 = _T_2699 ? _T_57556 : 16'h0; // @[Mux.scala 19:72:@28747.4]
  assign _T_57565 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5}; // @[Mux.scala 19:72:@28754.4]
  assign _T_57572 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13}; // @[Mux.scala 19:72:@28761.4]
  assign _T_57573 = {storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,_T_57565}; // @[Mux.scala 19:72:@28762.4]
  assign _T_57575 = _T_2700 ? _T_57573 : 16'h0; // @[Mux.scala 19:72:@28763.4]
  assign _T_57582 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6}; // @[Mux.scala 19:72:@28770.4]
  assign _T_57589 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14}; // @[Mux.scala 19:72:@28777.4]
  assign _T_57590 = {storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,storeAddrNotKnownFlags_6_14,_T_57582}; // @[Mux.scala 19:72:@28778.4]
  assign _T_57592 = _T_2701 ? _T_57590 : 16'h0; // @[Mux.scala 19:72:@28779.4]
  assign _T_57599 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7}; // @[Mux.scala 19:72:@28786.4]
  assign _T_57606 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15}; // @[Mux.scala 19:72:@28793.4]
  assign _T_57607 = {storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,storeAddrNotKnownFlags_6_15,_T_57599}; // @[Mux.scala 19:72:@28794.4]
  assign _T_57609 = _T_2702 ? _T_57607 : 16'h0; // @[Mux.scala 19:72:@28795.4]
  assign _T_57624 = {storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,storeAddrNotKnownFlags_6_0,_T_57487}; // @[Mux.scala 19:72:@28810.4]
  assign _T_57626 = _T_2703 ? _T_57624 : 16'h0; // @[Mux.scala 19:72:@28811.4]
  assign _T_57641 = {storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,storeAddrNotKnownFlags_6_1,_T_57504}; // @[Mux.scala 19:72:@28826.4]
  assign _T_57643 = _T_2704 ? _T_57641 : 16'h0; // @[Mux.scala 19:72:@28827.4]
  assign _T_57658 = {storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,storeAddrNotKnownFlags_6_2,_T_57521}; // @[Mux.scala 19:72:@28842.4]
  assign _T_57660 = _T_2705 ? _T_57658 : 16'h0; // @[Mux.scala 19:72:@28843.4]
  assign _T_57675 = {storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,storeAddrNotKnownFlags_6_3,_T_57538}; // @[Mux.scala 19:72:@28858.4]
  assign _T_57677 = _T_2706 ? _T_57675 : 16'h0; // @[Mux.scala 19:72:@28859.4]
  assign _T_57692 = {storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,storeAddrNotKnownFlags_6_4,_T_57555}; // @[Mux.scala 19:72:@28874.4]
  assign _T_57694 = _T_2707 ? _T_57692 : 16'h0; // @[Mux.scala 19:72:@28875.4]
  assign _T_57709 = {storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,storeAddrNotKnownFlags_6_5,_T_57572}; // @[Mux.scala 19:72:@28890.4]
  assign _T_57711 = _T_2708 ? _T_57709 : 16'h0; // @[Mux.scala 19:72:@28891.4]
  assign _T_57726 = {storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,storeAddrNotKnownFlags_6_6,_T_57589}; // @[Mux.scala 19:72:@28906.4]
  assign _T_57728 = _T_2709 ? _T_57726 : 16'h0; // @[Mux.scala 19:72:@28907.4]
  assign _T_57743 = {storeAddrNotKnownFlags_6_14,storeAddrNotKnownFlags_6_13,storeAddrNotKnownFlags_6_12,storeAddrNotKnownFlags_6_11,storeAddrNotKnownFlags_6_10,storeAddrNotKnownFlags_6_9,storeAddrNotKnownFlags_6_8,storeAddrNotKnownFlags_6_7,_T_57606}; // @[Mux.scala 19:72:@28922.4]
  assign _T_57745 = _T_2710 ? _T_57743 : 16'h0; // @[Mux.scala 19:72:@28923.4]
  assign _T_57746 = _T_57490 | _T_57507; // @[Mux.scala 19:72:@28924.4]
  assign _T_57747 = _T_57746 | _T_57524; // @[Mux.scala 19:72:@28925.4]
  assign _T_57748 = _T_57747 | _T_57541; // @[Mux.scala 19:72:@28926.4]
  assign _T_57749 = _T_57748 | _T_57558; // @[Mux.scala 19:72:@28927.4]
  assign _T_57750 = _T_57749 | _T_57575; // @[Mux.scala 19:72:@28928.4]
  assign _T_57751 = _T_57750 | _T_57592; // @[Mux.scala 19:72:@28929.4]
  assign _T_57752 = _T_57751 | _T_57609; // @[Mux.scala 19:72:@28930.4]
  assign _T_57753 = _T_57752 | _T_57626; // @[Mux.scala 19:72:@28931.4]
  assign _T_57754 = _T_57753 | _T_57643; // @[Mux.scala 19:72:@28932.4]
  assign _T_57755 = _T_57754 | _T_57660; // @[Mux.scala 19:72:@28933.4]
  assign _T_57756 = _T_57755 | _T_57677; // @[Mux.scala 19:72:@28934.4]
  assign _T_57757 = _T_57756 | _T_57694; // @[Mux.scala 19:72:@28935.4]
  assign _T_57758 = _T_57757 | _T_57711; // @[Mux.scala 19:72:@28936.4]
  assign _T_57759 = _T_57758 | _T_57728; // @[Mux.scala 19:72:@28937.4]
  assign _T_57760 = _T_57759 | _T_57745; // @[Mux.scala 19:72:@28938.4]
  assign _T_58338 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0}; // @[Mux.scala 19:72:@29288.4]
  assign _T_58345 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8}; // @[Mux.scala 19:72:@29295.4]
  assign _T_58346 = {storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,_T_58338}; // @[Mux.scala 19:72:@29296.4]
  assign _T_58348 = _T_2695 ? _T_58346 : 16'h0; // @[Mux.scala 19:72:@29297.4]
  assign _T_58355 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1}; // @[Mux.scala 19:72:@29304.4]
  assign _T_58362 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9}; // @[Mux.scala 19:72:@29311.4]
  assign _T_58363 = {storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,_T_58355}; // @[Mux.scala 19:72:@29312.4]
  assign _T_58365 = _T_2696 ? _T_58363 : 16'h0; // @[Mux.scala 19:72:@29313.4]
  assign _T_58372 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2}; // @[Mux.scala 19:72:@29320.4]
  assign _T_58379 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10}; // @[Mux.scala 19:72:@29327.4]
  assign _T_58380 = {storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,_T_58372}; // @[Mux.scala 19:72:@29328.4]
  assign _T_58382 = _T_2697 ? _T_58380 : 16'h0; // @[Mux.scala 19:72:@29329.4]
  assign _T_58389 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3}; // @[Mux.scala 19:72:@29336.4]
  assign _T_58396 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11}; // @[Mux.scala 19:72:@29343.4]
  assign _T_58397 = {storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,_T_58389}; // @[Mux.scala 19:72:@29344.4]
  assign _T_58399 = _T_2698 ? _T_58397 : 16'h0; // @[Mux.scala 19:72:@29345.4]
  assign _T_58406 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4}; // @[Mux.scala 19:72:@29352.4]
  assign _T_58413 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12}; // @[Mux.scala 19:72:@29359.4]
  assign _T_58414 = {storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,_T_58406}; // @[Mux.scala 19:72:@29360.4]
  assign _T_58416 = _T_2699 ? _T_58414 : 16'h0; // @[Mux.scala 19:72:@29361.4]
  assign _T_58423 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5}; // @[Mux.scala 19:72:@29368.4]
  assign _T_58430 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13}; // @[Mux.scala 19:72:@29375.4]
  assign _T_58431 = {storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,_T_58423}; // @[Mux.scala 19:72:@29376.4]
  assign _T_58433 = _T_2700 ? _T_58431 : 16'h0; // @[Mux.scala 19:72:@29377.4]
  assign _T_58440 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6}; // @[Mux.scala 19:72:@29384.4]
  assign _T_58447 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14}; // @[Mux.scala 19:72:@29391.4]
  assign _T_58448 = {storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,storeAddrNotKnownFlags_7_14,_T_58440}; // @[Mux.scala 19:72:@29392.4]
  assign _T_58450 = _T_2701 ? _T_58448 : 16'h0; // @[Mux.scala 19:72:@29393.4]
  assign _T_58457 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7}; // @[Mux.scala 19:72:@29400.4]
  assign _T_58464 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15}; // @[Mux.scala 19:72:@29407.4]
  assign _T_58465 = {storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,storeAddrNotKnownFlags_7_15,_T_58457}; // @[Mux.scala 19:72:@29408.4]
  assign _T_58467 = _T_2702 ? _T_58465 : 16'h0; // @[Mux.scala 19:72:@29409.4]
  assign _T_58482 = {storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,storeAddrNotKnownFlags_7_0,_T_58345}; // @[Mux.scala 19:72:@29424.4]
  assign _T_58484 = _T_2703 ? _T_58482 : 16'h0; // @[Mux.scala 19:72:@29425.4]
  assign _T_58499 = {storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,storeAddrNotKnownFlags_7_1,_T_58362}; // @[Mux.scala 19:72:@29440.4]
  assign _T_58501 = _T_2704 ? _T_58499 : 16'h0; // @[Mux.scala 19:72:@29441.4]
  assign _T_58516 = {storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,storeAddrNotKnownFlags_7_2,_T_58379}; // @[Mux.scala 19:72:@29456.4]
  assign _T_58518 = _T_2705 ? _T_58516 : 16'h0; // @[Mux.scala 19:72:@29457.4]
  assign _T_58533 = {storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,storeAddrNotKnownFlags_7_3,_T_58396}; // @[Mux.scala 19:72:@29472.4]
  assign _T_58535 = _T_2706 ? _T_58533 : 16'h0; // @[Mux.scala 19:72:@29473.4]
  assign _T_58550 = {storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,storeAddrNotKnownFlags_7_4,_T_58413}; // @[Mux.scala 19:72:@29488.4]
  assign _T_58552 = _T_2707 ? _T_58550 : 16'h0; // @[Mux.scala 19:72:@29489.4]
  assign _T_58567 = {storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,storeAddrNotKnownFlags_7_5,_T_58430}; // @[Mux.scala 19:72:@29504.4]
  assign _T_58569 = _T_2708 ? _T_58567 : 16'h0; // @[Mux.scala 19:72:@29505.4]
  assign _T_58584 = {storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,storeAddrNotKnownFlags_7_6,_T_58447}; // @[Mux.scala 19:72:@29520.4]
  assign _T_58586 = _T_2709 ? _T_58584 : 16'h0; // @[Mux.scala 19:72:@29521.4]
  assign _T_58601 = {storeAddrNotKnownFlags_7_14,storeAddrNotKnownFlags_7_13,storeAddrNotKnownFlags_7_12,storeAddrNotKnownFlags_7_11,storeAddrNotKnownFlags_7_10,storeAddrNotKnownFlags_7_9,storeAddrNotKnownFlags_7_8,storeAddrNotKnownFlags_7_7,_T_58464}; // @[Mux.scala 19:72:@29536.4]
  assign _T_58603 = _T_2710 ? _T_58601 : 16'h0; // @[Mux.scala 19:72:@29537.4]
  assign _T_58604 = _T_58348 | _T_58365; // @[Mux.scala 19:72:@29538.4]
  assign _T_58605 = _T_58604 | _T_58382; // @[Mux.scala 19:72:@29539.4]
  assign _T_58606 = _T_58605 | _T_58399; // @[Mux.scala 19:72:@29540.4]
  assign _T_58607 = _T_58606 | _T_58416; // @[Mux.scala 19:72:@29541.4]
  assign _T_58608 = _T_58607 | _T_58433; // @[Mux.scala 19:72:@29542.4]
  assign _T_58609 = _T_58608 | _T_58450; // @[Mux.scala 19:72:@29543.4]
  assign _T_58610 = _T_58609 | _T_58467; // @[Mux.scala 19:72:@29544.4]
  assign _T_58611 = _T_58610 | _T_58484; // @[Mux.scala 19:72:@29545.4]
  assign _T_58612 = _T_58611 | _T_58501; // @[Mux.scala 19:72:@29546.4]
  assign _T_58613 = _T_58612 | _T_58518; // @[Mux.scala 19:72:@29547.4]
  assign _T_58614 = _T_58613 | _T_58535; // @[Mux.scala 19:72:@29548.4]
  assign _T_58615 = _T_58614 | _T_58552; // @[Mux.scala 19:72:@29549.4]
  assign _T_58616 = _T_58615 | _T_58569; // @[Mux.scala 19:72:@29550.4]
  assign _T_58617 = _T_58616 | _T_58586; // @[Mux.scala 19:72:@29551.4]
  assign _T_58618 = _T_58617 | _T_58603; // @[Mux.scala 19:72:@29552.4]
  assign _T_59196 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0}; // @[Mux.scala 19:72:@29902.4]
  assign _T_59203 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8}; // @[Mux.scala 19:72:@29909.4]
  assign _T_59204 = {storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,_T_59196}; // @[Mux.scala 19:72:@29910.4]
  assign _T_59206 = _T_2695 ? _T_59204 : 16'h0; // @[Mux.scala 19:72:@29911.4]
  assign _T_59213 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1}; // @[Mux.scala 19:72:@29918.4]
  assign _T_59220 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9}; // @[Mux.scala 19:72:@29925.4]
  assign _T_59221 = {storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,_T_59213}; // @[Mux.scala 19:72:@29926.4]
  assign _T_59223 = _T_2696 ? _T_59221 : 16'h0; // @[Mux.scala 19:72:@29927.4]
  assign _T_59230 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2}; // @[Mux.scala 19:72:@29934.4]
  assign _T_59237 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10}; // @[Mux.scala 19:72:@29941.4]
  assign _T_59238 = {storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,_T_59230}; // @[Mux.scala 19:72:@29942.4]
  assign _T_59240 = _T_2697 ? _T_59238 : 16'h0; // @[Mux.scala 19:72:@29943.4]
  assign _T_59247 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3}; // @[Mux.scala 19:72:@29950.4]
  assign _T_59254 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11}; // @[Mux.scala 19:72:@29957.4]
  assign _T_59255 = {storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,_T_59247}; // @[Mux.scala 19:72:@29958.4]
  assign _T_59257 = _T_2698 ? _T_59255 : 16'h0; // @[Mux.scala 19:72:@29959.4]
  assign _T_59264 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4}; // @[Mux.scala 19:72:@29966.4]
  assign _T_59271 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12}; // @[Mux.scala 19:72:@29973.4]
  assign _T_59272 = {storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,_T_59264}; // @[Mux.scala 19:72:@29974.4]
  assign _T_59274 = _T_2699 ? _T_59272 : 16'h0; // @[Mux.scala 19:72:@29975.4]
  assign _T_59281 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5}; // @[Mux.scala 19:72:@29982.4]
  assign _T_59288 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13}; // @[Mux.scala 19:72:@29989.4]
  assign _T_59289 = {storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,_T_59281}; // @[Mux.scala 19:72:@29990.4]
  assign _T_59291 = _T_2700 ? _T_59289 : 16'h0; // @[Mux.scala 19:72:@29991.4]
  assign _T_59298 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6}; // @[Mux.scala 19:72:@29998.4]
  assign _T_59305 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14}; // @[Mux.scala 19:72:@30005.4]
  assign _T_59306 = {storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,storeAddrNotKnownFlags_8_14,_T_59298}; // @[Mux.scala 19:72:@30006.4]
  assign _T_59308 = _T_2701 ? _T_59306 : 16'h0; // @[Mux.scala 19:72:@30007.4]
  assign _T_59315 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7}; // @[Mux.scala 19:72:@30014.4]
  assign _T_59322 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15}; // @[Mux.scala 19:72:@30021.4]
  assign _T_59323 = {storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,storeAddrNotKnownFlags_8_15,_T_59315}; // @[Mux.scala 19:72:@30022.4]
  assign _T_59325 = _T_2702 ? _T_59323 : 16'h0; // @[Mux.scala 19:72:@30023.4]
  assign _T_59340 = {storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,storeAddrNotKnownFlags_8_0,_T_59203}; // @[Mux.scala 19:72:@30038.4]
  assign _T_59342 = _T_2703 ? _T_59340 : 16'h0; // @[Mux.scala 19:72:@30039.4]
  assign _T_59357 = {storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,storeAddrNotKnownFlags_8_1,_T_59220}; // @[Mux.scala 19:72:@30054.4]
  assign _T_59359 = _T_2704 ? _T_59357 : 16'h0; // @[Mux.scala 19:72:@30055.4]
  assign _T_59374 = {storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,storeAddrNotKnownFlags_8_2,_T_59237}; // @[Mux.scala 19:72:@30070.4]
  assign _T_59376 = _T_2705 ? _T_59374 : 16'h0; // @[Mux.scala 19:72:@30071.4]
  assign _T_59391 = {storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,storeAddrNotKnownFlags_8_3,_T_59254}; // @[Mux.scala 19:72:@30086.4]
  assign _T_59393 = _T_2706 ? _T_59391 : 16'h0; // @[Mux.scala 19:72:@30087.4]
  assign _T_59408 = {storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,storeAddrNotKnownFlags_8_4,_T_59271}; // @[Mux.scala 19:72:@30102.4]
  assign _T_59410 = _T_2707 ? _T_59408 : 16'h0; // @[Mux.scala 19:72:@30103.4]
  assign _T_59425 = {storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,storeAddrNotKnownFlags_8_5,_T_59288}; // @[Mux.scala 19:72:@30118.4]
  assign _T_59427 = _T_2708 ? _T_59425 : 16'h0; // @[Mux.scala 19:72:@30119.4]
  assign _T_59442 = {storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,storeAddrNotKnownFlags_8_6,_T_59305}; // @[Mux.scala 19:72:@30134.4]
  assign _T_59444 = _T_2709 ? _T_59442 : 16'h0; // @[Mux.scala 19:72:@30135.4]
  assign _T_59459 = {storeAddrNotKnownFlags_8_14,storeAddrNotKnownFlags_8_13,storeAddrNotKnownFlags_8_12,storeAddrNotKnownFlags_8_11,storeAddrNotKnownFlags_8_10,storeAddrNotKnownFlags_8_9,storeAddrNotKnownFlags_8_8,storeAddrNotKnownFlags_8_7,_T_59322}; // @[Mux.scala 19:72:@30150.4]
  assign _T_59461 = _T_2710 ? _T_59459 : 16'h0; // @[Mux.scala 19:72:@30151.4]
  assign _T_59462 = _T_59206 | _T_59223; // @[Mux.scala 19:72:@30152.4]
  assign _T_59463 = _T_59462 | _T_59240; // @[Mux.scala 19:72:@30153.4]
  assign _T_59464 = _T_59463 | _T_59257; // @[Mux.scala 19:72:@30154.4]
  assign _T_59465 = _T_59464 | _T_59274; // @[Mux.scala 19:72:@30155.4]
  assign _T_59466 = _T_59465 | _T_59291; // @[Mux.scala 19:72:@30156.4]
  assign _T_59467 = _T_59466 | _T_59308; // @[Mux.scala 19:72:@30157.4]
  assign _T_59468 = _T_59467 | _T_59325; // @[Mux.scala 19:72:@30158.4]
  assign _T_59469 = _T_59468 | _T_59342; // @[Mux.scala 19:72:@30159.4]
  assign _T_59470 = _T_59469 | _T_59359; // @[Mux.scala 19:72:@30160.4]
  assign _T_59471 = _T_59470 | _T_59376; // @[Mux.scala 19:72:@30161.4]
  assign _T_59472 = _T_59471 | _T_59393; // @[Mux.scala 19:72:@30162.4]
  assign _T_59473 = _T_59472 | _T_59410; // @[Mux.scala 19:72:@30163.4]
  assign _T_59474 = _T_59473 | _T_59427; // @[Mux.scala 19:72:@30164.4]
  assign _T_59475 = _T_59474 | _T_59444; // @[Mux.scala 19:72:@30165.4]
  assign _T_59476 = _T_59475 | _T_59461; // @[Mux.scala 19:72:@30166.4]
  assign _T_60054 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0}; // @[Mux.scala 19:72:@30516.4]
  assign _T_60061 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8}; // @[Mux.scala 19:72:@30523.4]
  assign _T_60062 = {storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,_T_60054}; // @[Mux.scala 19:72:@30524.4]
  assign _T_60064 = _T_2695 ? _T_60062 : 16'h0; // @[Mux.scala 19:72:@30525.4]
  assign _T_60071 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1}; // @[Mux.scala 19:72:@30532.4]
  assign _T_60078 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9}; // @[Mux.scala 19:72:@30539.4]
  assign _T_60079 = {storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,_T_60071}; // @[Mux.scala 19:72:@30540.4]
  assign _T_60081 = _T_2696 ? _T_60079 : 16'h0; // @[Mux.scala 19:72:@30541.4]
  assign _T_60088 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2}; // @[Mux.scala 19:72:@30548.4]
  assign _T_60095 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10}; // @[Mux.scala 19:72:@30555.4]
  assign _T_60096 = {storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,_T_60088}; // @[Mux.scala 19:72:@30556.4]
  assign _T_60098 = _T_2697 ? _T_60096 : 16'h0; // @[Mux.scala 19:72:@30557.4]
  assign _T_60105 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3}; // @[Mux.scala 19:72:@30564.4]
  assign _T_60112 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11}; // @[Mux.scala 19:72:@30571.4]
  assign _T_60113 = {storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,_T_60105}; // @[Mux.scala 19:72:@30572.4]
  assign _T_60115 = _T_2698 ? _T_60113 : 16'h0; // @[Mux.scala 19:72:@30573.4]
  assign _T_60122 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4}; // @[Mux.scala 19:72:@30580.4]
  assign _T_60129 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12}; // @[Mux.scala 19:72:@30587.4]
  assign _T_60130 = {storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,_T_60122}; // @[Mux.scala 19:72:@30588.4]
  assign _T_60132 = _T_2699 ? _T_60130 : 16'h0; // @[Mux.scala 19:72:@30589.4]
  assign _T_60139 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5}; // @[Mux.scala 19:72:@30596.4]
  assign _T_60146 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13}; // @[Mux.scala 19:72:@30603.4]
  assign _T_60147 = {storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,_T_60139}; // @[Mux.scala 19:72:@30604.4]
  assign _T_60149 = _T_2700 ? _T_60147 : 16'h0; // @[Mux.scala 19:72:@30605.4]
  assign _T_60156 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6}; // @[Mux.scala 19:72:@30612.4]
  assign _T_60163 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14}; // @[Mux.scala 19:72:@30619.4]
  assign _T_60164 = {storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,storeAddrNotKnownFlags_9_14,_T_60156}; // @[Mux.scala 19:72:@30620.4]
  assign _T_60166 = _T_2701 ? _T_60164 : 16'h0; // @[Mux.scala 19:72:@30621.4]
  assign _T_60173 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7}; // @[Mux.scala 19:72:@30628.4]
  assign _T_60180 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15}; // @[Mux.scala 19:72:@30635.4]
  assign _T_60181 = {storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,storeAddrNotKnownFlags_9_15,_T_60173}; // @[Mux.scala 19:72:@30636.4]
  assign _T_60183 = _T_2702 ? _T_60181 : 16'h0; // @[Mux.scala 19:72:@30637.4]
  assign _T_60198 = {storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,storeAddrNotKnownFlags_9_0,_T_60061}; // @[Mux.scala 19:72:@30652.4]
  assign _T_60200 = _T_2703 ? _T_60198 : 16'h0; // @[Mux.scala 19:72:@30653.4]
  assign _T_60215 = {storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,storeAddrNotKnownFlags_9_1,_T_60078}; // @[Mux.scala 19:72:@30668.4]
  assign _T_60217 = _T_2704 ? _T_60215 : 16'h0; // @[Mux.scala 19:72:@30669.4]
  assign _T_60232 = {storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,storeAddrNotKnownFlags_9_2,_T_60095}; // @[Mux.scala 19:72:@30684.4]
  assign _T_60234 = _T_2705 ? _T_60232 : 16'h0; // @[Mux.scala 19:72:@30685.4]
  assign _T_60249 = {storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,storeAddrNotKnownFlags_9_3,_T_60112}; // @[Mux.scala 19:72:@30700.4]
  assign _T_60251 = _T_2706 ? _T_60249 : 16'h0; // @[Mux.scala 19:72:@30701.4]
  assign _T_60266 = {storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,storeAddrNotKnownFlags_9_4,_T_60129}; // @[Mux.scala 19:72:@30716.4]
  assign _T_60268 = _T_2707 ? _T_60266 : 16'h0; // @[Mux.scala 19:72:@30717.4]
  assign _T_60283 = {storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,storeAddrNotKnownFlags_9_5,_T_60146}; // @[Mux.scala 19:72:@30732.4]
  assign _T_60285 = _T_2708 ? _T_60283 : 16'h0; // @[Mux.scala 19:72:@30733.4]
  assign _T_60300 = {storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,storeAddrNotKnownFlags_9_6,_T_60163}; // @[Mux.scala 19:72:@30748.4]
  assign _T_60302 = _T_2709 ? _T_60300 : 16'h0; // @[Mux.scala 19:72:@30749.4]
  assign _T_60317 = {storeAddrNotKnownFlags_9_14,storeAddrNotKnownFlags_9_13,storeAddrNotKnownFlags_9_12,storeAddrNotKnownFlags_9_11,storeAddrNotKnownFlags_9_10,storeAddrNotKnownFlags_9_9,storeAddrNotKnownFlags_9_8,storeAddrNotKnownFlags_9_7,_T_60180}; // @[Mux.scala 19:72:@30764.4]
  assign _T_60319 = _T_2710 ? _T_60317 : 16'h0; // @[Mux.scala 19:72:@30765.4]
  assign _T_60320 = _T_60064 | _T_60081; // @[Mux.scala 19:72:@30766.4]
  assign _T_60321 = _T_60320 | _T_60098; // @[Mux.scala 19:72:@30767.4]
  assign _T_60322 = _T_60321 | _T_60115; // @[Mux.scala 19:72:@30768.4]
  assign _T_60323 = _T_60322 | _T_60132; // @[Mux.scala 19:72:@30769.4]
  assign _T_60324 = _T_60323 | _T_60149; // @[Mux.scala 19:72:@30770.4]
  assign _T_60325 = _T_60324 | _T_60166; // @[Mux.scala 19:72:@30771.4]
  assign _T_60326 = _T_60325 | _T_60183; // @[Mux.scala 19:72:@30772.4]
  assign _T_60327 = _T_60326 | _T_60200; // @[Mux.scala 19:72:@30773.4]
  assign _T_60328 = _T_60327 | _T_60217; // @[Mux.scala 19:72:@30774.4]
  assign _T_60329 = _T_60328 | _T_60234; // @[Mux.scala 19:72:@30775.4]
  assign _T_60330 = _T_60329 | _T_60251; // @[Mux.scala 19:72:@30776.4]
  assign _T_60331 = _T_60330 | _T_60268; // @[Mux.scala 19:72:@30777.4]
  assign _T_60332 = _T_60331 | _T_60285; // @[Mux.scala 19:72:@30778.4]
  assign _T_60333 = _T_60332 | _T_60302; // @[Mux.scala 19:72:@30779.4]
  assign _T_60334 = _T_60333 | _T_60319; // @[Mux.scala 19:72:@30780.4]
  assign _T_60912 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0}; // @[Mux.scala 19:72:@31130.4]
  assign _T_60919 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8}; // @[Mux.scala 19:72:@31137.4]
  assign _T_60920 = {storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,_T_60912}; // @[Mux.scala 19:72:@31138.4]
  assign _T_60922 = _T_2695 ? _T_60920 : 16'h0; // @[Mux.scala 19:72:@31139.4]
  assign _T_60929 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1}; // @[Mux.scala 19:72:@31146.4]
  assign _T_60936 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9}; // @[Mux.scala 19:72:@31153.4]
  assign _T_60937 = {storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,_T_60929}; // @[Mux.scala 19:72:@31154.4]
  assign _T_60939 = _T_2696 ? _T_60937 : 16'h0; // @[Mux.scala 19:72:@31155.4]
  assign _T_60946 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2}; // @[Mux.scala 19:72:@31162.4]
  assign _T_60953 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10}; // @[Mux.scala 19:72:@31169.4]
  assign _T_60954 = {storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,_T_60946}; // @[Mux.scala 19:72:@31170.4]
  assign _T_60956 = _T_2697 ? _T_60954 : 16'h0; // @[Mux.scala 19:72:@31171.4]
  assign _T_60963 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3}; // @[Mux.scala 19:72:@31178.4]
  assign _T_60970 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11}; // @[Mux.scala 19:72:@31185.4]
  assign _T_60971 = {storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,_T_60963}; // @[Mux.scala 19:72:@31186.4]
  assign _T_60973 = _T_2698 ? _T_60971 : 16'h0; // @[Mux.scala 19:72:@31187.4]
  assign _T_60980 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4}; // @[Mux.scala 19:72:@31194.4]
  assign _T_60987 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12}; // @[Mux.scala 19:72:@31201.4]
  assign _T_60988 = {storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,_T_60980}; // @[Mux.scala 19:72:@31202.4]
  assign _T_60990 = _T_2699 ? _T_60988 : 16'h0; // @[Mux.scala 19:72:@31203.4]
  assign _T_60997 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5}; // @[Mux.scala 19:72:@31210.4]
  assign _T_61004 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13}; // @[Mux.scala 19:72:@31217.4]
  assign _T_61005 = {storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,_T_60997}; // @[Mux.scala 19:72:@31218.4]
  assign _T_61007 = _T_2700 ? _T_61005 : 16'h0; // @[Mux.scala 19:72:@31219.4]
  assign _T_61014 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6}; // @[Mux.scala 19:72:@31226.4]
  assign _T_61021 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14}; // @[Mux.scala 19:72:@31233.4]
  assign _T_61022 = {storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,storeAddrNotKnownFlags_10_14,_T_61014}; // @[Mux.scala 19:72:@31234.4]
  assign _T_61024 = _T_2701 ? _T_61022 : 16'h0; // @[Mux.scala 19:72:@31235.4]
  assign _T_61031 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7}; // @[Mux.scala 19:72:@31242.4]
  assign _T_61038 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15}; // @[Mux.scala 19:72:@31249.4]
  assign _T_61039 = {storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,storeAddrNotKnownFlags_10_15,_T_61031}; // @[Mux.scala 19:72:@31250.4]
  assign _T_61041 = _T_2702 ? _T_61039 : 16'h0; // @[Mux.scala 19:72:@31251.4]
  assign _T_61056 = {storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,storeAddrNotKnownFlags_10_0,_T_60919}; // @[Mux.scala 19:72:@31266.4]
  assign _T_61058 = _T_2703 ? _T_61056 : 16'h0; // @[Mux.scala 19:72:@31267.4]
  assign _T_61073 = {storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,storeAddrNotKnownFlags_10_1,_T_60936}; // @[Mux.scala 19:72:@31282.4]
  assign _T_61075 = _T_2704 ? _T_61073 : 16'h0; // @[Mux.scala 19:72:@31283.4]
  assign _T_61090 = {storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,storeAddrNotKnownFlags_10_2,_T_60953}; // @[Mux.scala 19:72:@31298.4]
  assign _T_61092 = _T_2705 ? _T_61090 : 16'h0; // @[Mux.scala 19:72:@31299.4]
  assign _T_61107 = {storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,storeAddrNotKnownFlags_10_3,_T_60970}; // @[Mux.scala 19:72:@31314.4]
  assign _T_61109 = _T_2706 ? _T_61107 : 16'h0; // @[Mux.scala 19:72:@31315.4]
  assign _T_61124 = {storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,storeAddrNotKnownFlags_10_4,_T_60987}; // @[Mux.scala 19:72:@31330.4]
  assign _T_61126 = _T_2707 ? _T_61124 : 16'h0; // @[Mux.scala 19:72:@31331.4]
  assign _T_61141 = {storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,storeAddrNotKnownFlags_10_5,_T_61004}; // @[Mux.scala 19:72:@31346.4]
  assign _T_61143 = _T_2708 ? _T_61141 : 16'h0; // @[Mux.scala 19:72:@31347.4]
  assign _T_61158 = {storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,storeAddrNotKnownFlags_10_6,_T_61021}; // @[Mux.scala 19:72:@31362.4]
  assign _T_61160 = _T_2709 ? _T_61158 : 16'h0; // @[Mux.scala 19:72:@31363.4]
  assign _T_61175 = {storeAddrNotKnownFlags_10_14,storeAddrNotKnownFlags_10_13,storeAddrNotKnownFlags_10_12,storeAddrNotKnownFlags_10_11,storeAddrNotKnownFlags_10_10,storeAddrNotKnownFlags_10_9,storeAddrNotKnownFlags_10_8,storeAddrNotKnownFlags_10_7,_T_61038}; // @[Mux.scala 19:72:@31378.4]
  assign _T_61177 = _T_2710 ? _T_61175 : 16'h0; // @[Mux.scala 19:72:@31379.4]
  assign _T_61178 = _T_60922 | _T_60939; // @[Mux.scala 19:72:@31380.4]
  assign _T_61179 = _T_61178 | _T_60956; // @[Mux.scala 19:72:@31381.4]
  assign _T_61180 = _T_61179 | _T_60973; // @[Mux.scala 19:72:@31382.4]
  assign _T_61181 = _T_61180 | _T_60990; // @[Mux.scala 19:72:@31383.4]
  assign _T_61182 = _T_61181 | _T_61007; // @[Mux.scala 19:72:@31384.4]
  assign _T_61183 = _T_61182 | _T_61024; // @[Mux.scala 19:72:@31385.4]
  assign _T_61184 = _T_61183 | _T_61041; // @[Mux.scala 19:72:@31386.4]
  assign _T_61185 = _T_61184 | _T_61058; // @[Mux.scala 19:72:@31387.4]
  assign _T_61186 = _T_61185 | _T_61075; // @[Mux.scala 19:72:@31388.4]
  assign _T_61187 = _T_61186 | _T_61092; // @[Mux.scala 19:72:@31389.4]
  assign _T_61188 = _T_61187 | _T_61109; // @[Mux.scala 19:72:@31390.4]
  assign _T_61189 = _T_61188 | _T_61126; // @[Mux.scala 19:72:@31391.4]
  assign _T_61190 = _T_61189 | _T_61143; // @[Mux.scala 19:72:@31392.4]
  assign _T_61191 = _T_61190 | _T_61160; // @[Mux.scala 19:72:@31393.4]
  assign _T_61192 = _T_61191 | _T_61177; // @[Mux.scala 19:72:@31394.4]
  assign _T_61770 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0}; // @[Mux.scala 19:72:@31744.4]
  assign _T_61777 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8}; // @[Mux.scala 19:72:@31751.4]
  assign _T_61778 = {storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,_T_61770}; // @[Mux.scala 19:72:@31752.4]
  assign _T_61780 = _T_2695 ? _T_61778 : 16'h0; // @[Mux.scala 19:72:@31753.4]
  assign _T_61787 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1}; // @[Mux.scala 19:72:@31760.4]
  assign _T_61794 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9}; // @[Mux.scala 19:72:@31767.4]
  assign _T_61795 = {storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,_T_61787}; // @[Mux.scala 19:72:@31768.4]
  assign _T_61797 = _T_2696 ? _T_61795 : 16'h0; // @[Mux.scala 19:72:@31769.4]
  assign _T_61804 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2}; // @[Mux.scala 19:72:@31776.4]
  assign _T_61811 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10}; // @[Mux.scala 19:72:@31783.4]
  assign _T_61812 = {storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,_T_61804}; // @[Mux.scala 19:72:@31784.4]
  assign _T_61814 = _T_2697 ? _T_61812 : 16'h0; // @[Mux.scala 19:72:@31785.4]
  assign _T_61821 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3}; // @[Mux.scala 19:72:@31792.4]
  assign _T_61828 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11}; // @[Mux.scala 19:72:@31799.4]
  assign _T_61829 = {storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,_T_61821}; // @[Mux.scala 19:72:@31800.4]
  assign _T_61831 = _T_2698 ? _T_61829 : 16'h0; // @[Mux.scala 19:72:@31801.4]
  assign _T_61838 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4}; // @[Mux.scala 19:72:@31808.4]
  assign _T_61845 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12}; // @[Mux.scala 19:72:@31815.4]
  assign _T_61846 = {storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,_T_61838}; // @[Mux.scala 19:72:@31816.4]
  assign _T_61848 = _T_2699 ? _T_61846 : 16'h0; // @[Mux.scala 19:72:@31817.4]
  assign _T_61855 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5}; // @[Mux.scala 19:72:@31824.4]
  assign _T_61862 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13}; // @[Mux.scala 19:72:@31831.4]
  assign _T_61863 = {storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,_T_61855}; // @[Mux.scala 19:72:@31832.4]
  assign _T_61865 = _T_2700 ? _T_61863 : 16'h0; // @[Mux.scala 19:72:@31833.4]
  assign _T_61872 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6}; // @[Mux.scala 19:72:@31840.4]
  assign _T_61879 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14}; // @[Mux.scala 19:72:@31847.4]
  assign _T_61880 = {storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,storeAddrNotKnownFlags_11_14,_T_61872}; // @[Mux.scala 19:72:@31848.4]
  assign _T_61882 = _T_2701 ? _T_61880 : 16'h0; // @[Mux.scala 19:72:@31849.4]
  assign _T_61889 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7}; // @[Mux.scala 19:72:@31856.4]
  assign _T_61896 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15}; // @[Mux.scala 19:72:@31863.4]
  assign _T_61897 = {storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,storeAddrNotKnownFlags_11_15,_T_61889}; // @[Mux.scala 19:72:@31864.4]
  assign _T_61899 = _T_2702 ? _T_61897 : 16'h0; // @[Mux.scala 19:72:@31865.4]
  assign _T_61914 = {storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,storeAddrNotKnownFlags_11_0,_T_61777}; // @[Mux.scala 19:72:@31880.4]
  assign _T_61916 = _T_2703 ? _T_61914 : 16'h0; // @[Mux.scala 19:72:@31881.4]
  assign _T_61931 = {storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,storeAddrNotKnownFlags_11_1,_T_61794}; // @[Mux.scala 19:72:@31896.4]
  assign _T_61933 = _T_2704 ? _T_61931 : 16'h0; // @[Mux.scala 19:72:@31897.4]
  assign _T_61948 = {storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,storeAddrNotKnownFlags_11_2,_T_61811}; // @[Mux.scala 19:72:@31912.4]
  assign _T_61950 = _T_2705 ? _T_61948 : 16'h0; // @[Mux.scala 19:72:@31913.4]
  assign _T_61965 = {storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,storeAddrNotKnownFlags_11_3,_T_61828}; // @[Mux.scala 19:72:@31928.4]
  assign _T_61967 = _T_2706 ? _T_61965 : 16'h0; // @[Mux.scala 19:72:@31929.4]
  assign _T_61982 = {storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,storeAddrNotKnownFlags_11_4,_T_61845}; // @[Mux.scala 19:72:@31944.4]
  assign _T_61984 = _T_2707 ? _T_61982 : 16'h0; // @[Mux.scala 19:72:@31945.4]
  assign _T_61999 = {storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,storeAddrNotKnownFlags_11_5,_T_61862}; // @[Mux.scala 19:72:@31960.4]
  assign _T_62001 = _T_2708 ? _T_61999 : 16'h0; // @[Mux.scala 19:72:@31961.4]
  assign _T_62016 = {storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,storeAddrNotKnownFlags_11_6,_T_61879}; // @[Mux.scala 19:72:@31976.4]
  assign _T_62018 = _T_2709 ? _T_62016 : 16'h0; // @[Mux.scala 19:72:@31977.4]
  assign _T_62033 = {storeAddrNotKnownFlags_11_14,storeAddrNotKnownFlags_11_13,storeAddrNotKnownFlags_11_12,storeAddrNotKnownFlags_11_11,storeAddrNotKnownFlags_11_10,storeAddrNotKnownFlags_11_9,storeAddrNotKnownFlags_11_8,storeAddrNotKnownFlags_11_7,_T_61896}; // @[Mux.scala 19:72:@31992.4]
  assign _T_62035 = _T_2710 ? _T_62033 : 16'h0; // @[Mux.scala 19:72:@31993.4]
  assign _T_62036 = _T_61780 | _T_61797; // @[Mux.scala 19:72:@31994.4]
  assign _T_62037 = _T_62036 | _T_61814; // @[Mux.scala 19:72:@31995.4]
  assign _T_62038 = _T_62037 | _T_61831; // @[Mux.scala 19:72:@31996.4]
  assign _T_62039 = _T_62038 | _T_61848; // @[Mux.scala 19:72:@31997.4]
  assign _T_62040 = _T_62039 | _T_61865; // @[Mux.scala 19:72:@31998.4]
  assign _T_62041 = _T_62040 | _T_61882; // @[Mux.scala 19:72:@31999.4]
  assign _T_62042 = _T_62041 | _T_61899; // @[Mux.scala 19:72:@32000.4]
  assign _T_62043 = _T_62042 | _T_61916; // @[Mux.scala 19:72:@32001.4]
  assign _T_62044 = _T_62043 | _T_61933; // @[Mux.scala 19:72:@32002.4]
  assign _T_62045 = _T_62044 | _T_61950; // @[Mux.scala 19:72:@32003.4]
  assign _T_62046 = _T_62045 | _T_61967; // @[Mux.scala 19:72:@32004.4]
  assign _T_62047 = _T_62046 | _T_61984; // @[Mux.scala 19:72:@32005.4]
  assign _T_62048 = _T_62047 | _T_62001; // @[Mux.scala 19:72:@32006.4]
  assign _T_62049 = _T_62048 | _T_62018; // @[Mux.scala 19:72:@32007.4]
  assign _T_62050 = _T_62049 | _T_62035; // @[Mux.scala 19:72:@32008.4]
  assign _T_62628 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0}; // @[Mux.scala 19:72:@32358.4]
  assign _T_62635 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8}; // @[Mux.scala 19:72:@32365.4]
  assign _T_62636 = {storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,_T_62628}; // @[Mux.scala 19:72:@32366.4]
  assign _T_62638 = _T_2695 ? _T_62636 : 16'h0; // @[Mux.scala 19:72:@32367.4]
  assign _T_62645 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1}; // @[Mux.scala 19:72:@32374.4]
  assign _T_62652 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9}; // @[Mux.scala 19:72:@32381.4]
  assign _T_62653 = {storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,_T_62645}; // @[Mux.scala 19:72:@32382.4]
  assign _T_62655 = _T_2696 ? _T_62653 : 16'h0; // @[Mux.scala 19:72:@32383.4]
  assign _T_62662 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2}; // @[Mux.scala 19:72:@32390.4]
  assign _T_62669 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10}; // @[Mux.scala 19:72:@32397.4]
  assign _T_62670 = {storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,_T_62662}; // @[Mux.scala 19:72:@32398.4]
  assign _T_62672 = _T_2697 ? _T_62670 : 16'h0; // @[Mux.scala 19:72:@32399.4]
  assign _T_62679 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3}; // @[Mux.scala 19:72:@32406.4]
  assign _T_62686 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11}; // @[Mux.scala 19:72:@32413.4]
  assign _T_62687 = {storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,_T_62679}; // @[Mux.scala 19:72:@32414.4]
  assign _T_62689 = _T_2698 ? _T_62687 : 16'h0; // @[Mux.scala 19:72:@32415.4]
  assign _T_62696 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4}; // @[Mux.scala 19:72:@32422.4]
  assign _T_62703 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12}; // @[Mux.scala 19:72:@32429.4]
  assign _T_62704 = {storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,_T_62696}; // @[Mux.scala 19:72:@32430.4]
  assign _T_62706 = _T_2699 ? _T_62704 : 16'h0; // @[Mux.scala 19:72:@32431.4]
  assign _T_62713 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5}; // @[Mux.scala 19:72:@32438.4]
  assign _T_62720 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13}; // @[Mux.scala 19:72:@32445.4]
  assign _T_62721 = {storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,_T_62713}; // @[Mux.scala 19:72:@32446.4]
  assign _T_62723 = _T_2700 ? _T_62721 : 16'h0; // @[Mux.scala 19:72:@32447.4]
  assign _T_62730 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6}; // @[Mux.scala 19:72:@32454.4]
  assign _T_62737 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14}; // @[Mux.scala 19:72:@32461.4]
  assign _T_62738 = {storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,storeAddrNotKnownFlags_12_14,_T_62730}; // @[Mux.scala 19:72:@32462.4]
  assign _T_62740 = _T_2701 ? _T_62738 : 16'h0; // @[Mux.scala 19:72:@32463.4]
  assign _T_62747 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7}; // @[Mux.scala 19:72:@32470.4]
  assign _T_62754 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15}; // @[Mux.scala 19:72:@32477.4]
  assign _T_62755 = {storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,storeAddrNotKnownFlags_12_15,_T_62747}; // @[Mux.scala 19:72:@32478.4]
  assign _T_62757 = _T_2702 ? _T_62755 : 16'h0; // @[Mux.scala 19:72:@32479.4]
  assign _T_62772 = {storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,storeAddrNotKnownFlags_12_0,_T_62635}; // @[Mux.scala 19:72:@32494.4]
  assign _T_62774 = _T_2703 ? _T_62772 : 16'h0; // @[Mux.scala 19:72:@32495.4]
  assign _T_62789 = {storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,storeAddrNotKnownFlags_12_1,_T_62652}; // @[Mux.scala 19:72:@32510.4]
  assign _T_62791 = _T_2704 ? _T_62789 : 16'h0; // @[Mux.scala 19:72:@32511.4]
  assign _T_62806 = {storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,storeAddrNotKnownFlags_12_2,_T_62669}; // @[Mux.scala 19:72:@32526.4]
  assign _T_62808 = _T_2705 ? _T_62806 : 16'h0; // @[Mux.scala 19:72:@32527.4]
  assign _T_62823 = {storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,storeAddrNotKnownFlags_12_3,_T_62686}; // @[Mux.scala 19:72:@32542.4]
  assign _T_62825 = _T_2706 ? _T_62823 : 16'h0; // @[Mux.scala 19:72:@32543.4]
  assign _T_62840 = {storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,storeAddrNotKnownFlags_12_4,_T_62703}; // @[Mux.scala 19:72:@32558.4]
  assign _T_62842 = _T_2707 ? _T_62840 : 16'h0; // @[Mux.scala 19:72:@32559.4]
  assign _T_62857 = {storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,storeAddrNotKnownFlags_12_5,_T_62720}; // @[Mux.scala 19:72:@32574.4]
  assign _T_62859 = _T_2708 ? _T_62857 : 16'h0; // @[Mux.scala 19:72:@32575.4]
  assign _T_62874 = {storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,storeAddrNotKnownFlags_12_6,_T_62737}; // @[Mux.scala 19:72:@32590.4]
  assign _T_62876 = _T_2709 ? _T_62874 : 16'h0; // @[Mux.scala 19:72:@32591.4]
  assign _T_62891 = {storeAddrNotKnownFlags_12_14,storeAddrNotKnownFlags_12_13,storeAddrNotKnownFlags_12_12,storeAddrNotKnownFlags_12_11,storeAddrNotKnownFlags_12_10,storeAddrNotKnownFlags_12_9,storeAddrNotKnownFlags_12_8,storeAddrNotKnownFlags_12_7,_T_62754}; // @[Mux.scala 19:72:@32606.4]
  assign _T_62893 = _T_2710 ? _T_62891 : 16'h0; // @[Mux.scala 19:72:@32607.4]
  assign _T_62894 = _T_62638 | _T_62655; // @[Mux.scala 19:72:@32608.4]
  assign _T_62895 = _T_62894 | _T_62672; // @[Mux.scala 19:72:@32609.4]
  assign _T_62896 = _T_62895 | _T_62689; // @[Mux.scala 19:72:@32610.4]
  assign _T_62897 = _T_62896 | _T_62706; // @[Mux.scala 19:72:@32611.4]
  assign _T_62898 = _T_62897 | _T_62723; // @[Mux.scala 19:72:@32612.4]
  assign _T_62899 = _T_62898 | _T_62740; // @[Mux.scala 19:72:@32613.4]
  assign _T_62900 = _T_62899 | _T_62757; // @[Mux.scala 19:72:@32614.4]
  assign _T_62901 = _T_62900 | _T_62774; // @[Mux.scala 19:72:@32615.4]
  assign _T_62902 = _T_62901 | _T_62791; // @[Mux.scala 19:72:@32616.4]
  assign _T_62903 = _T_62902 | _T_62808; // @[Mux.scala 19:72:@32617.4]
  assign _T_62904 = _T_62903 | _T_62825; // @[Mux.scala 19:72:@32618.4]
  assign _T_62905 = _T_62904 | _T_62842; // @[Mux.scala 19:72:@32619.4]
  assign _T_62906 = _T_62905 | _T_62859; // @[Mux.scala 19:72:@32620.4]
  assign _T_62907 = _T_62906 | _T_62876; // @[Mux.scala 19:72:@32621.4]
  assign _T_62908 = _T_62907 | _T_62893; // @[Mux.scala 19:72:@32622.4]
  assign _T_63486 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0}; // @[Mux.scala 19:72:@32972.4]
  assign _T_63493 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8}; // @[Mux.scala 19:72:@32979.4]
  assign _T_63494 = {storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,_T_63486}; // @[Mux.scala 19:72:@32980.4]
  assign _T_63496 = _T_2695 ? _T_63494 : 16'h0; // @[Mux.scala 19:72:@32981.4]
  assign _T_63503 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1}; // @[Mux.scala 19:72:@32988.4]
  assign _T_63510 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9}; // @[Mux.scala 19:72:@32995.4]
  assign _T_63511 = {storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,_T_63503}; // @[Mux.scala 19:72:@32996.4]
  assign _T_63513 = _T_2696 ? _T_63511 : 16'h0; // @[Mux.scala 19:72:@32997.4]
  assign _T_63520 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2}; // @[Mux.scala 19:72:@33004.4]
  assign _T_63527 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10}; // @[Mux.scala 19:72:@33011.4]
  assign _T_63528 = {storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,_T_63520}; // @[Mux.scala 19:72:@33012.4]
  assign _T_63530 = _T_2697 ? _T_63528 : 16'h0; // @[Mux.scala 19:72:@33013.4]
  assign _T_63537 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3}; // @[Mux.scala 19:72:@33020.4]
  assign _T_63544 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11}; // @[Mux.scala 19:72:@33027.4]
  assign _T_63545 = {storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,_T_63537}; // @[Mux.scala 19:72:@33028.4]
  assign _T_63547 = _T_2698 ? _T_63545 : 16'h0; // @[Mux.scala 19:72:@33029.4]
  assign _T_63554 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4}; // @[Mux.scala 19:72:@33036.4]
  assign _T_63561 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12}; // @[Mux.scala 19:72:@33043.4]
  assign _T_63562 = {storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,_T_63554}; // @[Mux.scala 19:72:@33044.4]
  assign _T_63564 = _T_2699 ? _T_63562 : 16'h0; // @[Mux.scala 19:72:@33045.4]
  assign _T_63571 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5}; // @[Mux.scala 19:72:@33052.4]
  assign _T_63578 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13}; // @[Mux.scala 19:72:@33059.4]
  assign _T_63579 = {storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,_T_63571}; // @[Mux.scala 19:72:@33060.4]
  assign _T_63581 = _T_2700 ? _T_63579 : 16'h0; // @[Mux.scala 19:72:@33061.4]
  assign _T_63588 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6}; // @[Mux.scala 19:72:@33068.4]
  assign _T_63595 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14}; // @[Mux.scala 19:72:@33075.4]
  assign _T_63596 = {storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,storeAddrNotKnownFlags_13_14,_T_63588}; // @[Mux.scala 19:72:@33076.4]
  assign _T_63598 = _T_2701 ? _T_63596 : 16'h0; // @[Mux.scala 19:72:@33077.4]
  assign _T_63605 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7}; // @[Mux.scala 19:72:@33084.4]
  assign _T_63612 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15}; // @[Mux.scala 19:72:@33091.4]
  assign _T_63613 = {storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,storeAddrNotKnownFlags_13_15,_T_63605}; // @[Mux.scala 19:72:@33092.4]
  assign _T_63615 = _T_2702 ? _T_63613 : 16'h0; // @[Mux.scala 19:72:@33093.4]
  assign _T_63630 = {storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,storeAddrNotKnownFlags_13_0,_T_63493}; // @[Mux.scala 19:72:@33108.4]
  assign _T_63632 = _T_2703 ? _T_63630 : 16'h0; // @[Mux.scala 19:72:@33109.4]
  assign _T_63647 = {storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,storeAddrNotKnownFlags_13_1,_T_63510}; // @[Mux.scala 19:72:@33124.4]
  assign _T_63649 = _T_2704 ? _T_63647 : 16'h0; // @[Mux.scala 19:72:@33125.4]
  assign _T_63664 = {storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,storeAddrNotKnownFlags_13_2,_T_63527}; // @[Mux.scala 19:72:@33140.4]
  assign _T_63666 = _T_2705 ? _T_63664 : 16'h0; // @[Mux.scala 19:72:@33141.4]
  assign _T_63681 = {storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,storeAddrNotKnownFlags_13_3,_T_63544}; // @[Mux.scala 19:72:@33156.4]
  assign _T_63683 = _T_2706 ? _T_63681 : 16'h0; // @[Mux.scala 19:72:@33157.4]
  assign _T_63698 = {storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,storeAddrNotKnownFlags_13_4,_T_63561}; // @[Mux.scala 19:72:@33172.4]
  assign _T_63700 = _T_2707 ? _T_63698 : 16'h0; // @[Mux.scala 19:72:@33173.4]
  assign _T_63715 = {storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,storeAddrNotKnownFlags_13_5,_T_63578}; // @[Mux.scala 19:72:@33188.4]
  assign _T_63717 = _T_2708 ? _T_63715 : 16'h0; // @[Mux.scala 19:72:@33189.4]
  assign _T_63732 = {storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,storeAddrNotKnownFlags_13_6,_T_63595}; // @[Mux.scala 19:72:@33204.4]
  assign _T_63734 = _T_2709 ? _T_63732 : 16'h0; // @[Mux.scala 19:72:@33205.4]
  assign _T_63749 = {storeAddrNotKnownFlags_13_14,storeAddrNotKnownFlags_13_13,storeAddrNotKnownFlags_13_12,storeAddrNotKnownFlags_13_11,storeAddrNotKnownFlags_13_10,storeAddrNotKnownFlags_13_9,storeAddrNotKnownFlags_13_8,storeAddrNotKnownFlags_13_7,_T_63612}; // @[Mux.scala 19:72:@33220.4]
  assign _T_63751 = _T_2710 ? _T_63749 : 16'h0; // @[Mux.scala 19:72:@33221.4]
  assign _T_63752 = _T_63496 | _T_63513; // @[Mux.scala 19:72:@33222.4]
  assign _T_63753 = _T_63752 | _T_63530; // @[Mux.scala 19:72:@33223.4]
  assign _T_63754 = _T_63753 | _T_63547; // @[Mux.scala 19:72:@33224.4]
  assign _T_63755 = _T_63754 | _T_63564; // @[Mux.scala 19:72:@33225.4]
  assign _T_63756 = _T_63755 | _T_63581; // @[Mux.scala 19:72:@33226.4]
  assign _T_63757 = _T_63756 | _T_63598; // @[Mux.scala 19:72:@33227.4]
  assign _T_63758 = _T_63757 | _T_63615; // @[Mux.scala 19:72:@33228.4]
  assign _T_63759 = _T_63758 | _T_63632; // @[Mux.scala 19:72:@33229.4]
  assign _T_63760 = _T_63759 | _T_63649; // @[Mux.scala 19:72:@33230.4]
  assign _T_63761 = _T_63760 | _T_63666; // @[Mux.scala 19:72:@33231.4]
  assign _T_63762 = _T_63761 | _T_63683; // @[Mux.scala 19:72:@33232.4]
  assign _T_63763 = _T_63762 | _T_63700; // @[Mux.scala 19:72:@33233.4]
  assign _T_63764 = _T_63763 | _T_63717; // @[Mux.scala 19:72:@33234.4]
  assign _T_63765 = _T_63764 | _T_63734; // @[Mux.scala 19:72:@33235.4]
  assign _T_63766 = _T_63765 | _T_63751; // @[Mux.scala 19:72:@33236.4]
  assign _T_64344 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0}; // @[Mux.scala 19:72:@33586.4]
  assign _T_64351 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8}; // @[Mux.scala 19:72:@33593.4]
  assign _T_64352 = {storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,_T_64344}; // @[Mux.scala 19:72:@33594.4]
  assign _T_64354 = _T_2695 ? _T_64352 : 16'h0; // @[Mux.scala 19:72:@33595.4]
  assign _T_64361 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1}; // @[Mux.scala 19:72:@33602.4]
  assign _T_64368 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9}; // @[Mux.scala 19:72:@33609.4]
  assign _T_64369 = {storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,_T_64361}; // @[Mux.scala 19:72:@33610.4]
  assign _T_64371 = _T_2696 ? _T_64369 : 16'h0; // @[Mux.scala 19:72:@33611.4]
  assign _T_64378 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2}; // @[Mux.scala 19:72:@33618.4]
  assign _T_64385 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10}; // @[Mux.scala 19:72:@33625.4]
  assign _T_64386 = {storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,_T_64378}; // @[Mux.scala 19:72:@33626.4]
  assign _T_64388 = _T_2697 ? _T_64386 : 16'h0; // @[Mux.scala 19:72:@33627.4]
  assign _T_64395 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3}; // @[Mux.scala 19:72:@33634.4]
  assign _T_64402 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11}; // @[Mux.scala 19:72:@33641.4]
  assign _T_64403 = {storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,_T_64395}; // @[Mux.scala 19:72:@33642.4]
  assign _T_64405 = _T_2698 ? _T_64403 : 16'h0; // @[Mux.scala 19:72:@33643.4]
  assign _T_64412 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4}; // @[Mux.scala 19:72:@33650.4]
  assign _T_64419 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12}; // @[Mux.scala 19:72:@33657.4]
  assign _T_64420 = {storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,_T_64412}; // @[Mux.scala 19:72:@33658.4]
  assign _T_64422 = _T_2699 ? _T_64420 : 16'h0; // @[Mux.scala 19:72:@33659.4]
  assign _T_64429 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5}; // @[Mux.scala 19:72:@33666.4]
  assign _T_64436 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13}; // @[Mux.scala 19:72:@33673.4]
  assign _T_64437 = {storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,_T_64429}; // @[Mux.scala 19:72:@33674.4]
  assign _T_64439 = _T_2700 ? _T_64437 : 16'h0; // @[Mux.scala 19:72:@33675.4]
  assign _T_64446 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6}; // @[Mux.scala 19:72:@33682.4]
  assign _T_64453 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14}; // @[Mux.scala 19:72:@33689.4]
  assign _T_64454 = {storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,storeAddrNotKnownFlags_14_14,_T_64446}; // @[Mux.scala 19:72:@33690.4]
  assign _T_64456 = _T_2701 ? _T_64454 : 16'h0; // @[Mux.scala 19:72:@33691.4]
  assign _T_64463 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7}; // @[Mux.scala 19:72:@33698.4]
  assign _T_64470 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15}; // @[Mux.scala 19:72:@33705.4]
  assign _T_64471 = {storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,storeAddrNotKnownFlags_14_15,_T_64463}; // @[Mux.scala 19:72:@33706.4]
  assign _T_64473 = _T_2702 ? _T_64471 : 16'h0; // @[Mux.scala 19:72:@33707.4]
  assign _T_64488 = {storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,storeAddrNotKnownFlags_14_0,_T_64351}; // @[Mux.scala 19:72:@33722.4]
  assign _T_64490 = _T_2703 ? _T_64488 : 16'h0; // @[Mux.scala 19:72:@33723.4]
  assign _T_64505 = {storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,storeAddrNotKnownFlags_14_1,_T_64368}; // @[Mux.scala 19:72:@33738.4]
  assign _T_64507 = _T_2704 ? _T_64505 : 16'h0; // @[Mux.scala 19:72:@33739.4]
  assign _T_64522 = {storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,storeAddrNotKnownFlags_14_2,_T_64385}; // @[Mux.scala 19:72:@33754.4]
  assign _T_64524 = _T_2705 ? _T_64522 : 16'h0; // @[Mux.scala 19:72:@33755.4]
  assign _T_64539 = {storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,storeAddrNotKnownFlags_14_3,_T_64402}; // @[Mux.scala 19:72:@33770.4]
  assign _T_64541 = _T_2706 ? _T_64539 : 16'h0; // @[Mux.scala 19:72:@33771.4]
  assign _T_64556 = {storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,storeAddrNotKnownFlags_14_4,_T_64419}; // @[Mux.scala 19:72:@33786.4]
  assign _T_64558 = _T_2707 ? _T_64556 : 16'h0; // @[Mux.scala 19:72:@33787.4]
  assign _T_64573 = {storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,storeAddrNotKnownFlags_14_5,_T_64436}; // @[Mux.scala 19:72:@33802.4]
  assign _T_64575 = _T_2708 ? _T_64573 : 16'h0; // @[Mux.scala 19:72:@33803.4]
  assign _T_64590 = {storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,storeAddrNotKnownFlags_14_6,_T_64453}; // @[Mux.scala 19:72:@33818.4]
  assign _T_64592 = _T_2709 ? _T_64590 : 16'h0; // @[Mux.scala 19:72:@33819.4]
  assign _T_64607 = {storeAddrNotKnownFlags_14_14,storeAddrNotKnownFlags_14_13,storeAddrNotKnownFlags_14_12,storeAddrNotKnownFlags_14_11,storeAddrNotKnownFlags_14_10,storeAddrNotKnownFlags_14_9,storeAddrNotKnownFlags_14_8,storeAddrNotKnownFlags_14_7,_T_64470}; // @[Mux.scala 19:72:@33834.4]
  assign _T_64609 = _T_2710 ? _T_64607 : 16'h0; // @[Mux.scala 19:72:@33835.4]
  assign _T_64610 = _T_64354 | _T_64371; // @[Mux.scala 19:72:@33836.4]
  assign _T_64611 = _T_64610 | _T_64388; // @[Mux.scala 19:72:@33837.4]
  assign _T_64612 = _T_64611 | _T_64405; // @[Mux.scala 19:72:@33838.4]
  assign _T_64613 = _T_64612 | _T_64422; // @[Mux.scala 19:72:@33839.4]
  assign _T_64614 = _T_64613 | _T_64439; // @[Mux.scala 19:72:@33840.4]
  assign _T_64615 = _T_64614 | _T_64456; // @[Mux.scala 19:72:@33841.4]
  assign _T_64616 = _T_64615 | _T_64473; // @[Mux.scala 19:72:@33842.4]
  assign _T_64617 = _T_64616 | _T_64490; // @[Mux.scala 19:72:@33843.4]
  assign _T_64618 = _T_64617 | _T_64507; // @[Mux.scala 19:72:@33844.4]
  assign _T_64619 = _T_64618 | _T_64524; // @[Mux.scala 19:72:@33845.4]
  assign _T_64620 = _T_64619 | _T_64541; // @[Mux.scala 19:72:@33846.4]
  assign _T_64621 = _T_64620 | _T_64558; // @[Mux.scala 19:72:@33847.4]
  assign _T_64622 = _T_64621 | _T_64575; // @[Mux.scala 19:72:@33848.4]
  assign _T_64623 = _T_64622 | _T_64592; // @[Mux.scala 19:72:@33849.4]
  assign _T_64624 = _T_64623 | _T_64609; // @[Mux.scala 19:72:@33850.4]
  assign _T_65202 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0}; // @[Mux.scala 19:72:@34200.4]
  assign _T_65209 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8}; // @[Mux.scala 19:72:@34207.4]
  assign _T_65210 = {storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,_T_65202}; // @[Mux.scala 19:72:@34208.4]
  assign _T_65212 = _T_2695 ? _T_65210 : 16'h0; // @[Mux.scala 19:72:@34209.4]
  assign _T_65219 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1}; // @[Mux.scala 19:72:@34216.4]
  assign _T_65226 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9}; // @[Mux.scala 19:72:@34223.4]
  assign _T_65227 = {storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,_T_65219}; // @[Mux.scala 19:72:@34224.4]
  assign _T_65229 = _T_2696 ? _T_65227 : 16'h0; // @[Mux.scala 19:72:@34225.4]
  assign _T_65236 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2}; // @[Mux.scala 19:72:@34232.4]
  assign _T_65243 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10}; // @[Mux.scala 19:72:@34239.4]
  assign _T_65244 = {storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,_T_65236}; // @[Mux.scala 19:72:@34240.4]
  assign _T_65246 = _T_2697 ? _T_65244 : 16'h0; // @[Mux.scala 19:72:@34241.4]
  assign _T_65253 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3}; // @[Mux.scala 19:72:@34248.4]
  assign _T_65260 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11}; // @[Mux.scala 19:72:@34255.4]
  assign _T_65261 = {storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,_T_65253}; // @[Mux.scala 19:72:@34256.4]
  assign _T_65263 = _T_2698 ? _T_65261 : 16'h0; // @[Mux.scala 19:72:@34257.4]
  assign _T_65270 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4}; // @[Mux.scala 19:72:@34264.4]
  assign _T_65277 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12}; // @[Mux.scala 19:72:@34271.4]
  assign _T_65278 = {storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,_T_65270}; // @[Mux.scala 19:72:@34272.4]
  assign _T_65280 = _T_2699 ? _T_65278 : 16'h0; // @[Mux.scala 19:72:@34273.4]
  assign _T_65287 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5}; // @[Mux.scala 19:72:@34280.4]
  assign _T_65294 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13}; // @[Mux.scala 19:72:@34287.4]
  assign _T_65295 = {storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,_T_65287}; // @[Mux.scala 19:72:@34288.4]
  assign _T_65297 = _T_2700 ? _T_65295 : 16'h0; // @[Mux.scala 19:72:@34289.4]
  assign _T_65304 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6}; // @[Mux.scala 19:72:@34296.4]
  assign _T_65311 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14}; // @[Mux.scala 19:72:@34303.4]
  assign _T_65312 = {storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,storeAddrNotKnownFlags_15_14,_T_65304}; // @[Mux.scala 19:72:@34304.4]
  assign _T_65314 = _T_2701 ? _T_65312 : 16'h0; // @[Mux.scala 19:72:@34305.4]
  assign _T_65321 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7}; // @[Mux.scala 19:72:@34312.4]
  assign _T_65328 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15}; // @[Mux.scala 19:72:@34319.4]
  assign _T_65329 = {storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,storeAddrNotKnownFlags_15_15,_T_65321}; // @[Mux.scala 19:72:@34320.4]
  assign _T_65331 = _T_2702 ? _T_65329 : 16'h0; // @[Mux.scala 19:72:@34321.4]
  assign _T_65346 = {storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,storeAddrNotKnownFlags_15_0,_T_65209}; // @[Mux.scala 19:72:@34336.4]
  assign _T_65348 = _T_2703 ? _T_65346 : 16'h0; // @[Mux.scala 19:72:@34337.4]
  assign _T_65363 = {storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,storeAddrNotKnownFlags_15_1,_T_65226}; // @[Mux.scala 19:72:@34352.4]
  assign _T_65365 = _T_2704 ? _T_65363 : 16'h0; // @[Mux.scala 19:72:@34353.4]
  assign _T_65380 = {storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,storeAddrNotKnownFlags_15_2,_T_65243}; // @[Mux.scala 19:72:@34368.4]
  assign _T_65382 = _T_2705 ? _T_65380 : 16'h0; // @[Mux.scala 19:72:@34369.4]
  assign _T_65397 = {storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,storeAddrNotKnownFlags_15_3,_T_65260}; // @[Mux.scala 19:72:@34384.4]
  assign _T_65399 = _T_2706 ? _T_65397 : 16'h0; // @[Mux.scala 19:72:@34385.4]
  assign _T_65414 = {storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,storeAddrNotKnownFlags_15_4,_T_65277}; // @[Mux.scala 19:72:@34400.4]
  assign _T_65416 = _T_2707 ? _T_65414 : 16'h0; // @[Mux.scala 19:72:@34401.4]
  assign _T_65431 = {storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,storeAddrNotKnownFlags_15_5,_T_65294}; // @[Mux.scala 19:72:@34416.4]
  assign _T_65433 = _T_2708 ? _T_65431 : 16'h0; // @[Mux.scala 19:72:@34417.4]
  assign _T_65448 = {storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,storeAddrNotKnownFlags_15_6,_T_65311}; // @[Mux.scala 19:72:@34432.4]
  assign _T_65450 = _T_2709 ? _T_65448 : 16'h0; // @[Mux.scala 19:72:@34433.4]
  assign _T_65465 = {storeAddrNotKnownFlags_15_14,storeAddrNotKnownFlags_15_13,storeAddrNotKnownFlags_15_12,storeAddrNotKnownFlags_15_11,storeAddrNotKnownFlags_15_10,storeAddrNotKnownFlags_15_9,storeAddrNotKnownFlags_15_8,storeAddrNotKnownFlags_15_7,_T_65328}; // @[Mux.scala 19:72:@34448.4]
  assign _T_65467 = _T_2710 ? _T_65465 : 16'h0; // @[Mux.scala 19:72:@34449.4]
  assign _T_65468 = _T_65212 | _T_65229; // @[Mux.scala 19:72:@34450.4]
  assign _T_65469 = _T_65468 | _T_65246; // @[Mux.scala 19:72:@34451.4]
  assign _T_65470 = _T_65469 | _T_65263; // @[Mux.scala 19:72:@34452.4]
  assign _T_65471 = _T_65470 | _T_65280; // @[Mux.scala 19:72:@34453.4]
  assign _T_65472 = _T_65471 | _T_65297; // @[Mux.scala 19:72:@34454.4]
  assign _T_65473 = _T_65472 | _T_65314; // @[Mux.scala 19:72:@34455.4]
  assign _T_65474 = _T_65473 | _T_65331; // @[Mux.scala 19:72:@34456.4]
  assign _T_65475 = _T_65474 | _T_65348; // @[Mux.scala 19:72:@34457.4]
  assign _T_65476 = _T_65475 | _T_65365; // @[Mux.scala 19:72:@34458.4]
  assign _T_65477 = _T_65476 | _T_65382; // @[Mux.scala 19:72:@34459.4]
  assign _T_65478 = _T_65477 | _T_65399; // @[Mux.scala 19:72:@34460.4]
  assign _T_65479 = _T_65478 | _T_65416; // @[Mux.scala 19:72:@34461.4]
  assign _T_65480 = _T_65479 | _T_65433; // @[Mux.scala 19:72:@34462.4]
  assign _T_65481 = _T_65480 | _T_65450; // @[Mux.scala 19:72:@34463.4]
  assign _T_65482 = _T_65481 | _T_65467; // @[Mux.scala 19:72:@34464.4]
  assign _T_88274 = conflictPReg_0_2 ? 2'h2 : {{1'd0}, conflictPReg_0_1}; // @[AxiLoadQueue.scala 191:60:@35137.4]
  assign _T_88275 = conflictPReg_0_3 ? 2'h3 : _T_88274; // @[AxiLoadQueue.scala 191:60:@35138.4]
  assign _T_88276 = conflictPReg_0_4 ? 3'h4 : {{1'd0}, _T_88275}; // @[AxiLoadQueue.scala 191:60:@35139.4]
  assign _T_88277 = conflictPReg_0_5 ? 3'h5 : _T_88276; // @[AxiLoadQueue.scala 191:60:@35140.4]
  assign _T_88278 = conflictPReg_0_6 ? 3'h6 : _T_88277; // @[AxiLoadQueue.scala 191:60:@35141.4]
  assign _T_88279 = conflictPReg_0_7 ? 3'h7 : _T_88278; // @[AxiLoadQueue.scala 191:60:@35142.4]
  assign _T_88280 = conflictPReg_0_8 ? 4'h8 : {{1'd0}, _T_88279}; // @[AxiLoadQueue.scala 191:60:@35143.4]
  assign _T_88281 = conflictPReg_0_9 ? 4'h9 : _T_88280; // @[AxiLoadQueue.scala 191:60:@35144.4]
  assign _T_88282 = conflictPReg_0_10 ? 4'ha : _T_88281; // @[AxiLoadQueue.scala 191:60:@35145.4]
  assign _T_88283 = conflictPReg_0_11 ? 4'hb : _T_88282; // @[AxiLoadQueue.scala 191:60:@35146.4]
  assign _T_88284 = conflictPReg_0_12 ? 4'hc : _T_88283; // @[AxiLoadQueue.scala 191:60:@35147.4]
  assign _T_88285 = conflictPReg_0_13 ? 4'hd : _T_88284; // @[AxiLoadQueue.scala 191:60:@35148.4]
  assign _T_88286 = conflictPReg_0_14 ? 4'he : _T_88285; // @[AxiLoadQueue.scala 191:60:@35149.4]
  assign _T_88287 = conflictPReg_0_15 ? 4'hf : _T_88286; // @[AxiLoadQueue.scala 191:60:@35150.4]
  assign _T_88290 = conflictPReg_0_0 | conflictPReg_0_1; // @[AxiLoadQueue.scala 192:43:@35152.4]
  assign _T_88291 = _T_88290 | conflictPReg_0_2; // @[AxiLoadQueue.scala 192:43:@35153.4]
  assign _T_88292 = _T_88291 | conflictPReg_0_3; // @[AxiLoadQueue.scala 192:43:@35154.4]
  assign _T_88293 = _T_88292 | conflictPReg_0_4; // @[AxiLoadQueue.scala 192:43:@35155.4]
  assign _T_88294 = _T_88293 | conflictPReg_0_5; // @[AxiLoadQueue.scala 192:43:@35156.4]
  assign _T_88295 = _T_88294 | conflictPReg_0_6; // @[AxiLoadQueue.scala 192:43:@35157.4]
  assign _T_88296 = _T_88295 | conflictPReg_0_7; // @[AxiLoadQueue.scala 192:43:@35158.4]
  assign _T_88297 = _T_88296 | conflictPReg_0_8; // @[AxiLoadQueue.scala 192:43:@35159.4]
  assign _T_88298 = _T_88297 | conflictPReg_0_9; // @[AxiLoadQueue.scala 192:43:@35160.4]
  assign _T_88299 = _T_88298 | conflictPReg_0_10; // @[AxiLoadQueue.scala 192:43:@35161.4]
  assign _T_88300 = _T_88299 | conflictPReg_0_11; // @[AxiLoadQueue.scala 192:43:@35162.4]
  assign _T_88301 = _T_88300 | conflictPReg_0_12; // @[AxiLoadQueue.scala 192:43:@35163.4]
  assign _T_88302 = _T_88301 | conflictPReg_0_13; // @[AxiLoadQueue.scala 192:43:@35164.4]
  assign _T_88303 = _T_88302 | conflictPReg_0_14; // @[AxiLoadQueue.scala 192:43:@35165.4]
  assign _T_88304 = _T_88303 | conflictPReg_0_15; // @[AxiLoadQueue.scala 192:43:@35166.4]
  assign _GEN_864 = 4'h0 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_865 = 4'h1 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_866 = 4'h2 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_867 = 4'h3 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_868 = 4'h4 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_869 = 4'h5 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_870 = 4'h6 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_871 = 4'h7 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_872 = 4'h8 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_873 = 4'h9 == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_874 = 4'ha == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_875 = 4'hb == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_876 = 4'hc == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_877 = 4'hd == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_878 = 4'he == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_879 = 4'hf == _T_88287; // @[AxiLoadQueue.scala 193:43:@35168.6]
  assign _GEN_881 = 4'h1 == _T_88287 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_882 = 4'h2 == _T_88287 ? shiftedStoreDataKnownPReg_2 : _GEN_881; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_883 = 4'h3 == _T_88287 ? shiftedStoreDataKnownPReg_3 : _GEN_882; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_884 = 4'h4 == _T_88287 ? shiftedStoreDataKnownPReg_4 : _GEN_883; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_885 = 4'h5 == _T_88287 ? shiftedStoreDataKnownPReg_5 : _GEN_884; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_886 = 4'h6 == _T_88287 ? shiftedStoreDataKnownPReg_6 : _GEN_885; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_887 = 4'h7 == _T_88287 ? shiftedStoreDataKnownPReg_7 : _GEN_886; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_888 = 4'h8 == _T_88287 ? shiftedStoreDataKnownPReg_8 : _GEN_887; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_889 = 4'h9 == _T_88287 ? shiftedStoreDataKnownPReg_9 : _GEN_888; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_890 = 4'ha == _T_88287 ? shiftedStoreDataKnownPReg_10 : _GEN_889; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_891 = 4'hb == _T_88287 ? shiftedStoreDataKnownPReg_11 : _GEN_890; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_892 = 4'hc == _T_88287 ? shiftedStoreDataKnownPReg_12 : _GEN_891; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_893 = 4'hd == _T_88287 ? shiftedStoreDataKnownPReg_13 : _GEN_892; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_894 = 4'he == _T_88287 ? shiftedStoreDataKnownPReg_14 : _GEN_893; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_895 = 4'hf == _T_88287 ? shiftedStoreDataKnownPReg_15 : _GEN_894; // @[AxiLoadQueue.scala 194:31:@35169.6]
  assign _GEN_897 = 4'h1 == _T_88287 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_898 = 4'h2 == _T_88287 ? shiftedStoreDataQPreg_2 : _GEN_897; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_899 = 4'h3 == _T_88287 ? shiftedStoreDataQPreg_3 : _GEN_898; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_900 = 4'h4 == _T_88287 ? shiftedStoreDataQPreg_4 : _GEN_899; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_901 = 4'h5 == _T_88287 ? shiftedStoreDataQPreg_5 : _GEN_900; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_902 = 4'h6 == _T_88287 ? shiftedStoreDataQPreg_6 : _GEN_901; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_903 = 4'h7 == _T_88287 ? shiftedStoreDataQPreg_7 : _GEN_902; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_904 = 4'h8 == _T_88287 ? shiftedStoreDataQPreg_8 : _GEN_903; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_905 = 4'h9 == _T_88287 ? shiftedStoreDataQPreg_9 : _GEN_904; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_906 = 4'ha == _T_88287 ? shiftedStoreDataQPreg_10 : _GEN_905; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_907 = 4'hb == _T_88287 ? shiftedStoreDataQPreg_11 : _GEN_906; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_908 = 4'hc == _T_88287 ? shiftedStoreDataQPreg_12 : _GEN_907; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_909 = 4'hd == _T_88287 ? shiftedStoreDataQPreg_13 : _GEN_908; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_910 = 4'he == _T_88287 ? shiftedStoreDataQPreg_14 : _GEN_909; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign _GEN_911 = 4'hf == _T_88287 ? shiftedStoreDataQPreg_15 : _GEN_910; // @[AxiLoadQueue.scala 195:31:@35170.6]
  assign lastConflict_0_0 = _T_88304 ? _GEN_864 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_1 = _T_88304 ? _GEN_865 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_2 = _T_88304 ? _GEN_866 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_3 = _T_88304 ? _GEN_867 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_4 = _T_88304 ? _GEN_868 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_5 = _T_88304 ? _GEN_869 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_6 = _T_88304 ? _GEN_870 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_7 = _T_88304 ? _GEN_871 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_8 = _T_88304 ? _GEN_872 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_9 = _T_88304 ? _GEN_873 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_10 = _T_88304 ? _GEN_874 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_11 = _T_88304 ? _GEN_875 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_12 = _T_88304 ? _GEN_876 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_13 = _T_88304 ? _GEN_877 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_14 = _T_88304 ? _GEN_878 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign lastConflict_0_15 = _T_88304 ? _GEN_879 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign canBypass_0 = _T_88304 ? _GEN_895 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign bypassVal_0 = _T_88304 ? _GEN_911 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35167.4]
  assign _T_88410 = conflictPReg_1_2 ? 2'h2 : {{1'd0}, conflictPReg_1_1}; // @[AxiLoadQueue.scala 191:60:@35224.4]
  assign _T_88411 = conflictPReg_1_3 ? 2'h3 : _T_88410; // @[AxiLoadQueue.scala 191:60:@35225.4]
  assign _T_88412 = conflictPReg_1_4 ? 3'h4 : {{1'd0}, _T_88411}; // @[AxiLoadQueue.scala 191:60:@35226.4]
  assign _T_88413 = conflictPReg_1_5 ? 3'h5 : _T_88412; // @[AxiLoadQueue.scala 191:60:@35227.4]
  assign _T_88414 = conflictPReg_1_6 ? 3'h6 : _T_88413; // @[AxiLoadQueue.scala 191:60:@35228.4]
  assign _T_88415 = conflictPReg_1_7 ? 3'h7 : _T_88414; // @[AxiLoadQueue.scala 191:60:@35229.4]
  assign _T_88416 = conflictPReg_1_8 ? 4'h8 : {{1'd0}, _T_88415}; // @[AxiLoadQueue.scala 191:60:@35230.4]
  assign _T_88417 = conflictPReg_1_9 ? 4'h9 : _T_88416; // @[AxiLoadQueue.scala 191:60:@35231.4]
  assign _T_88418 = conflictPReg_1_10 ? 4'ha : _T_88417; // @[AxiLoadQueue.scala 191:60:@35232.4]
  assign _T_88419 = conflictPReg_1_11 ? 4'hb : _T_88418; // @[AxiLoadQueue.scala 191:60:@35233.4]
  assign _T_88420 = conflictPReg_1_12 ? 4'hc : _T_88419; // @[AxiLoadQueue.scala 191:60:@35234.4]
  assign _T_88421 = conflictPReg_1_13 ? 4'hd : _T_88420; // @[AxiLoadQueue.scala 191:60:@35235.4]
  assign _T_88422 = conflictPReg_1_14 ? 4'he : _T_88421; // @[AxiLoadQueue.scala 191:60:@35236.4]
  assign _T_88423 = conflictPReg_1_15 ? 4'hf : _T_88422; // @[AxiLoadQueue.scala 191:60:@35237.4]
  assign _T_88426 = conflictPReg_1_0 | conflictPReg_1_1; // @[AxiLoadQueue.scala 192:43:@35239.4]
  assign _T_88427 = _T_88426 | conflictPReg_1_2; // @[AxiLoadQueue.scala 192:43:@35240.4]
  assign _T_88428 = _T_88427 | conflictPReg_1_3; // @[AxiLoadQueue.scala 192:43:@35241.4]
  assign _T_88429 = _T_88428 | conflictPReg_1_4; // @[AxiLoadQueue.scala 192:43:@35242.4]
  assign _T_88430 = _T_88429 | conflictPReg_1_5; // @[AxiLoadQueue.scala 192:43:@35243.4]
  assign _T_88431 = _T_88430 | conflictPReg_1_6; // @[AxiLoadQueue.scala 192:43:@35244.4]
  assign _T_88432 = _T_88431 | conflictPReg_1_7; // @[AxiLoadQueue.scala 192:43:@35245.4]
  assign _T_88433 = _T_88432 | conflictPReg_1_8; // @[AxiLoadQueue.scala 192:43:@35246.4]
  assign _T_88434 = _T_88433 | conflictPReg_1_9; // @[AxiLoadQueue.scala 192:43:@35247.4]
  assign _T_88435 = _T_88434 | conflictPReg_1_10; // @[AxiLoadQueue.scala 192:43:@35248.4]
  assign _T_88436 = _T_88435 | conflictPReg_1_11; // @[AxiLoadQueue.scala 192:43:@35249.4]
  assign _T_88437 = _T_88436 | conflictPReg_1_12; // @[AxiLoadQueue.scala 192:43:@35250.4]
  assign _T_88438 = _T_88437 | conflictPReg_1_13; // @[AxiLoadQueue.scala 192:43:@35251.4]
  assign _T_88439 = _T_88438 | conflictPReg_1_14; // @[AxiLoadQueue.scala 192:43:@35252.4]
  assign _T_88440 = _T_88439 | conflictPReg_1_15; // @[AxiLoadQueue.scala 192:43:@35253.4]
  assign _GEN_930 = 4'h0 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_931 = 4'h1 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_932 = 4'h2 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_933 = 4'h3 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_934 = 4'h4 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_935 = 4'h5 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_936 = 4'h6 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_937 = 4'h7 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_938 = 4'h8 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_939 = 4'h9 == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_940 = 4'ha == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_941 = 4'hb == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_942 = 4'hc == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_943 = 4'hd == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_944 = 4'he == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_945 = 4'hf == _T_88423; // @[AxiLoadQueue.scala 193:43:@35255.6]
  assign _GEN_947 = 4'h1 == _T_88423 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_948 = 4'h2 == _T_88423 ? shiftedStoreDataKnownPReg_2 : _GEN_947; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_949 = 4'h3 == _T_88423 ? shiftedStoreDataKnownPReg_3 : _GEN_948; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_950 = 4'h4 == _T_88423 ? shiftedStoreDataKnownPReg_4 : _GEN_949; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_951 = 4'h5 == _T_88423 ? shiftedStoreDataKnownPReg_5 : _GEN_950; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_952 = 4'h6 == _T_88423 ? shiftedStoreDataKnownPReg_6 : _GEN_951; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_953 = 4'h7 == _T_88423 ? shiftedStoreDataKnownPReg_7 : _GEN_952; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_954 = 4'h8 == _T_88423 ? shiftedStoreDataKnownPReg_8 : _GEN_953; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_955 = 4'h9 == _T_88423 ? shiftedStoreDataKnownPReg_9 : _GEN_954; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_956 = 4'ha == _T_88423 ? shiftedStoreDataKnownPReg_10 : _GEN_955; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_957 = 4'hb == _T_88423 ? shiftedStoreDataKnownPReg_11 : _GEN_956; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_958 = 4'hc == _T_88423 ? shiftedStoreDataKnownPReg_12 : _GEN_957; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_959 = 4'hd == _T_88423 ? shiftedStoreDataKnownPReg_13 : _GEN_958; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_960 = 4'he == _T_88423 ? shiftedStoreDataKnownPReg_14 : _GEN_959; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_961 = 4'hf == _T_88423 ? shiftedStoreDataKnownPReg_15 : _GEN_960; // @[AxiLoadQueue.scala 194:31:@35256.6]
  assign _GEN_963 = 4'h1 == _T_88423 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_964 = 4'h2 == _T_88423 ? shiftedStoreDataQPreg_2 : _GEN_963; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_965 = 4'h3 == _T_88423 ? shiftedStoreDataQPreg_3 : _GEN_964; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_966 = 4'h4 == _T_88423 ? shiftedStoreDataQPreg_4 : _GEN_965; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_967 = 4'h5 == _T_88423 ? shiftedStoreDataQPreg_5 : _GEN_966; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_968 = 4'h6 == _T_88423 ? shiftedStoreDataQPreg_6 : _GEN_967; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_969 = 4'h7 == _T_88423 ? shiftedStoreDataQPreg_7 : _GEN_968; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_970 = 4'h8 == _T_88423 ? shiftedStoreDataQPreg_8 : _GEN_969; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_971 = 4'h9 == _T_88423 ? shiftedStoreDataQPreg_9 : _GEN_970; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_972 = 4'ha == _T_88423 ? shiftedStoreDataQPreg_10 : _GEN_971; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_973 = 4'hb == _T_88423 ? shiftedStoreDataQPreg_11 : _GEN_972; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_974 = 4'hc == _T_88423 ? shiftedStoreDataQPreg_12 : _GEN_973; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_975 = 4'hd == _T_88423 ? shiftedStoreDataQPreg_13 : _GEN_974; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_976 = 4'he == _T_88423 ? shiftedStoreDataQPreg_14 : _GEN_975; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign _GEN_977 = 4'hf == _T_88423 ? shiftedStoreDataQPreg_15 : _GEN_976; // @[AxiLoadQueue.scala 195:31:@35257.6]
  assign lastConflict_1_0 = _T_88440 ? _GEN_930 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_1 = _T_88440 ? _GEN_931 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_2 = _T_88440 ? _GEN_932 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_3 = _T_88440 ? _GEN_933 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_4 = _T_88440 ? _GEN_934 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_5 = _T_88440 ? _GEN_935 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_6 = _T_88440 ? _GEN_936 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_7 = _T_88440 ? _GEN_937 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_8 = _T_88440 ? _GEN_938 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_9 = _T_88440 ? _GEN_939 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_10 = _T_88440 ? _GEN_940 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_11 = _T_88440 ? _GEN_941 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_12 = _T_88440 ? _GEN_942 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_13 = _T_88440 ? _GEN_943 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_14 = _T_88440 ? _GEN_944 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign lastConflict_1_15 = _T_88440 ? _GEN_945 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign canBypass_1 = _T_88440 ? _GEN_961 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign bypassVal_1 = _T_88440 ? _GEN_977 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35254.4]
  assign _T_88546 = conflictPReg_2_2 ? 2'h2 : {{1'd0}, conflictPReg_2_1}; // @[AxiLoadQueue.scala 191:60:@35311.4]
  assign _T_88547 = conflictPReg_2_3 ? 2'h3 : _T_88546; // @[AxiLoadQueue.scala 191:60:@35312.4]
  assign _T_88548 = conflictPReg_2_4 ? 3'h4 : {{1'd0}, _T_88547}; // @[AxiLoadQueue.scala 191:60:@35313.4]
  assign _T_88549 = conflictPReg_2_5 ? 3'h5 : _T_88548; // @[AxiLoadQueue.scala 191:60:@35314.4]
  assign _T_88550 = conflictPReg_2_6 ? 3'h6 : _T_88549; // @[AxiLoadQueue.scala 191:60:@35315.4]
  assign _T_88551 = conflictPReg_2_7 ? 3'h7 : _T_88550; // @[AxiLoadQueue.scala 191:60:@35316.4]
  assign _T_88552 = conflictPReg_2_8 ? 4'h8 : {{1'd0}, _T_88551}; // @[AxiLoadQueue.scala 191:60:@35317.4]
  assign _T_88553 = conflictPReg_2_9 ? 4'h9 : _T_88552; // @[AxiLoadQueue.scala 191:60:@35318.4]
  assign _T_88554 = conflictPReg_2_10 ? 4'ha : _T_88553; // @[AxiLoadQueue.scala 191:60:@35319.4]
  assign _T_88555 = conflictPReg_2_11 ? 4'hb : _T_88554; // @[AxiLoadQueue.scala 191:60:@35320.4]
  assign _T_88556 = conflictPReg_2_12 ? 4'hc : _T_88555; // @[AxiLoadQueue.scala 191:60:@35321.4]
  assign _T_88557 = conflictPReg_2_13 ? 4'hd : _T_88556; // @[AxiLoadQueue.scala 191:60:@35322.4]
  assign _T_88558 = conflictPReg_2_14 ? 4'he : _T_88557; // @[AxiLoadQueue.scala 191:60:@35323.4]
  assign _T_88559 = conflictPReg_2_15 ? 4'hf : _T_88558; // @[AxiLoadQueue.scala 191:60:@35324.4]
  assign _T_88562 = conflictPReg_2_0 | conflictPReg_2_1; // @[AxiLoadQueue.scala 192:43:@35326.4]
  assign _T_88563 = _T_88562 | conflictPReg_2_2; // @[AxiLoadQueue.scala 192:43:@35327.4]
  assign _T_88564 = _T_88563 | conflictPReg_2_3; // @[AxiLoadQueue.scala 192:43:@35328.4]
  assign _T_88565 = _T_88564 | conflictPReg_2_4; // @[AxiLoadQueue.scala 192:43:@35329.4]
  assign _T_88566 = _T_88565 | conflictPReg_2_5; // @[AxiLoadQueue.scala 192:43:@35330.4]
  assign _T_88567 = _T_88566 | conflictPReg_2_6; // @[AxiLoadQueue.scala 192:43:@35331.4]
  assign _T_88568 = _T_88567 | conflictPReg_2_7; // @[AxiLoadQueue.scala 192:43:@35332.4]
  assign _T_88569 = _T_88568 | conflictPReg_2_8; // @[AxiLoadQueue.scala 192:43:@35333.4]
  assign _T_88570 = _T_88569 | conflictPReg_2_9; // @[AxiLoadQueue.scala 192:43:@35334.4]
  assign _T_88571 = _T_88570 | conflictPReg_2_10; // @[AxiLoadQueue.scala 192:43:@35335.4]
  assign _T_88572 = _T_88571 | conflictPReg_2_11; // @[AxiLoadQueue.scala 192:43:@35336.4]
  assign _T_88573 = _T_88572 | conflictPReg_2_12; // @[AxiLoadQueue.scala 192:43:@35337.4]
  assign _T_88574 = _T_88573 | conflictPReg_2_13; // @[AxiLoadQueue.scala 192:43:@35338.4]
  assign _T_88575 = _T_88574 | conflictPReg_2_14; // @[AxiLoadQueue.scala 192:43:@35339.4]
  assign _T_88576 = _T_88575 | conflictPReg_2_15; // @[AxiLoadQueue.scala 192:43:@35340.4]
  assign _GEN_996 = 4'h0 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_997 = 4'h1 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_998 = 4'h2 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_999 = 4'h3 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1000 = 4'h4 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1001 = 4'h5 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1002 = 4'h6 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1003 = 4'h7 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1004 = 4'h8 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1005 = 4'h9 == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1006 = 4'ha == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1007 = 4'hb == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1008 = 4'hc == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1009 = 4'hd == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1010 = 4'he == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1011 = 4'hf == _T_88559; // @[AxiLoadQueue.scala 193:43:@35342.6]
  assign _GEN_1013 = 4'h1 == _T_88559 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1014 = 4'h2 == _T_88559 ? shiftedStoreDataKnownPReg_2 : _GEN_1013; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1015 = 4'h3 == _T_88559 ? shiftedStoreDataKnownPReg_3 : _GEN_1014; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1016 = 4'h4 == _T_88559 ? shiftedStoreDataKnownPReg_4 : _GEN_1015; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1017 = 4'h5 == _T_88559 ? shiftedStoreDataKnownPReg_5 : _GEN_1016; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1018 = 4'h6 == _T_88559 ? shiftedStoreDataKnownPReg_6 : _GEN_1017; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1019 = 4'h7 == _T_88559 ? shiftedStoreDataKnownPReg_7 : _GEN_1018; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1020 = 4'h8 == _T_88559 ? shiftedStoreDataKnownPReg_8 : _GEN_1019; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1021 = 4'h9 == _T_88559 ? shiftedStoreDataKnownPReg_9 : _GEN_1020; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1022 = 4'ha == _T_88559 ? shiftedStoreDataKnownPReg_10 : _GEN_1021; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1023 = 4'hb == _T_88559 ? shiftedStoreDataKnownPReg_11 : _GEN_1022; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1024 = 4'hc == _T_88559 ? shiftedStoreDataKnownPReg_12 : _GEN_1023; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1025 = 4'hd == _T_88559 ? shiftedStoreDataKnownPReg_13 : _GEN_1024; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1026 = 4'he == _T_88559 ? shiftedStoreDataKnownPReg_14 : _GEN_1025; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1027 = 4'hf == _T_88559 ? shiftedStoreDataKnownPReg_15 : _GEN_1026; // @[AxiLoadQueue.scala 194:31:@35343.6]
  assign _GEN_1029 = 4'h1 == _T_88559 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1030 = 4'h2 == _T_88559 ? shiftedStoreDataQPreg_2 : _GEN_1029; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1031 = 4'h3 == _T_88559 ? shiftedStoreDataQPreg_3 : _GEN_1030; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1032 = 4'h4 == _T_88559 ? shiftedStoreDataQPreg_4 : _GEN_1031; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1033 = 4'h5 == _T_88559 ? shiftedStoreDataQPreg_5 : _GEN_1032; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1034 = 4'h6 == _T_88559 ? shiftedStoreDataQPreg_6 : _GEN_1033; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1035 = 4'h7 == _T_88559 ? shiftedStoreDataQPreg_7 : _GEN_1034; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1036 = 4'h8 == _T_88559 ? shiftedStoreDataQPreg_8 : _GEN_1035; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1037 = 4'h9 == _T_88559 ? shiftedStoreDataQPreg_9 : _GEN_1036; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1038 = 4'ha == _T_88559 ? shiftedStoreDataQPreg_10 : _GEN_1037; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1039 = 4'hb == _T_88559 ? shiftedStoreDataQPreg_11 : _GEN_1038; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1040 = 4'hc == _T_88559 ? shiftedStoreDataQPreg_12 : _GEN_1039; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1041 = 4'hd == _T_88559 ? shiftedStoreDataQPreg_13 : _GEN_1040; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1042 = 4'he == _T_88559 ? shiftedStoreDataQPreg_14 : _GEN_1041; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign _GEN_1043 = 4'hf == _T_88559 ? shiftedStoreDataQPreg_15 : _GEN_1042; // @[AxiLoadQueue.scala 195:31:@35344.6]
  assign lastConflict_2_0 = _T_88576 ? _GEN_996 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_1 = _T_88576 ? _GEN_997 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_2 = _T_88576 ? _GEN_998 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_3 = _T_88576 ? _GEN_999 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_4 = _T_88576 ? _GEN_1000 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_5 = _T_88576 ? _GEN_1001 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_6 = _T_88576 ? _GEN_1002 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_7 = _T_88576 ? _GEN_1003 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_8 = _T_88576 ? _GEN_1004 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_9 = _T_88576 ? _GEN_1005 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_10 = _T_88576 ? _GEN_1006 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_11 = _T_88576 ? _GEN_1007 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_12 = _T_88576 ? _GEN_1008 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_13 = _T_88576 ? _GEN_1009 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_14 = _T_88576 ? _GEN_1010 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign lastConflict_2_15 = _T_88576 ? _GEN_1011 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign canBypass_2 = _T_88576 ? _GEN_1027 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign bypassVal_2 = _T_88576 ? _GEN_1043 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35341.4]
  assign _T_88682 = conflictPReg_3_2 ? 2'h2 : {{1'd0}, conflictPReg_3_1}; // @[AxiLoadQueue.scala 191:60:@35398.4]
  assign _T_88683 = conflictPReg_3_3 ? 2'h3 : _T_88682; // @[AxiLoadQueue.scala 191:60:@35399.4]
  assign _T_88684 = conflictPReg_3_4 ? 3'h4 : {{1'd0}, _T_88683}; // @[AxiLoadQueue.scala 191:60:@35400.4]
  assign _T_88685 = conflictPReg_3_5 ? 3'h5 : _T_88684; // @[AxiLoadQueue.scala 191:60:@35401.4]
  assign _T_88686 = conflictPReg_3_6 ? 3'h6 : _T_88685; // @[AxiLoadQueue.scala 191:60:@35402.4]
  assign _T_88687 = conflictPReg_3_7 ? 3'h7 : _T_88686; // @[AxiLoadQueue.scala 191:60:@35403.4]
  assign _T_88688 = conflictPReg_3_8 ? 4'h8 : {{1'd0}, _T_88687}; // @[AxiLoadQueue.scala 191:60:@35404.4]
  assign _T_88689 = conflictPReg_3_9 ? 4'h9 : _T_88688; // @[AxiLoadQueue.scala 191:60:@35405.4]
  assign _T_88690 = conflictPReg_3_10 ? 4'ha : _T_88689; // @[AxiLoadQueue.scala 191:60:@35406.4]
  assign _T_88691 = conflictPReg_3_11 ? 4'hb : _T_88690; // @[AxiLoadQueue.scala 191:60:@35407.4]
  assign _T_88692 = conflictPReg_3_12 ? 4'hc : _T_88691; // @[AxiLoadQueue.scala 191:60:@35408.4]
  assign _T_88693 = conflictPReg_3_13 ? 4'hd : _T_88692; // @[AxiLoadQueue.scala 191:60:@35409.4]
  assign _T_88694 = conflictPReg_3_14 ? 4'he : _T_88693; // @[AxiLoadQueue.scala 191:60:@35410.4]
  assign _T_88695 = conflictPReg_3_15 ? 4'hf : _T_88694; // @[AxiLoadQueue.scala 191:60:@35411.4]
  assign _T_88698 = conflictPReg_3_0 | conflictPReg_3_1; // @[AxiLoadQueue.scala 192:43:@35413.4]
  assign _T_88699 = _T_88698 | conflictPReg_3_2; // @[AxiLoadQueue.scala 192:43:@35414.4]
  assign _T_88700 = _T_88699 | conflictPReg_3_3; // @[AxiLoadQueue.scala 192:43:@35415.4]
  assign _T_88701 = _T_88700 | conflictPReg_3_4; // @[AxiLoadQueue.scala 192:43:@35416.4]
  assign _T_88702 = _T_88701 | conflictPReg_3_5; // @[AxiLoadQueue.scala 192:43:@35417.4]
  assign _T_88703 = _T_88702 | conflictPReg_3_6; // @[AxiLoadQueue.scala 192:43:@35418.4]
  assign _T_88704 = _T_88703 | conflictPReg_3_7; // @[AxiLoadQueue.scala 192:43:@35419.4]
  assign _T_88705 = _T_88704 | conflictPReg_3_8; // @[AxiLoadQueue.scala 192:43:@35420.4]
  assign _T_88706 = _T_88705 | conflictPReg_3_9; // @[AxiLoadQueue.scala 192:43:@35421.4]
  assign _T_88707 = _T_88706 | conflictPReg_3_10; // @[AxiLoadQueue.scala 192:43:@35422.4]
  assign _T_88708 = _T_88707 | conflictPReg_3_11; // @[AxiLoadQueue.scala 192:43:@35423.4]
  assign _T_88709 = _T_88708 | conflictPReg_3_12; // @[AxiLoadQueue.scala 192:43:@35424.4]
  assign _T_88710 = _T_88709 | conflictPReg_3_13; // @[AxiLoadQueue.scala 192:43:@35425.4]
  assign _T_88711 = _T_88710 | conflictPReg_3_14; // @[AxiLoadQueue.scala 192:43:@35426.4]
  assign _T_88712 = _T_88711 | conflictPReg_3_15; // @[AxiLoadQueue.scala 192:43:@35427.4]
  assign _GEN_1062 = 4'h0 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1063 = 4'h1 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1064 = 4'h2 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1065 = 4'h3 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1066 = 4'h4 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1067 = 4'h5 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1068 = 4'h6 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1069 = 4'h7 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1070 = 4'h8 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1071 = 4'h9 == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1072 = 4'ha == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1073 = 4'hb == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1074 = 4'hc == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1075 = 4'hd == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1076 = 4'he == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1077 = 4'hf == _T_88695; // @[AxiLoadQueue.scala 193:43:@35429.6]
  assign _GEN_1079 = 4'h1 == _T_88695 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1080 = 4'h2 == _T_88695 ? shiftedStoreDataKnownPReg_2 : _GEN_1079; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1081 = 4'h3 == _T_88695 ? shiftedStoreDataKnownPReg_3 : _GEN_1080; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1082 = 4'h4 == _T_88695 ? shiftedStoreDataKnownPReg_4 : _GEN_1081; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1083 = 4'h5 == _T_88695 ? shiftedStoreDataKnownPReg_5 : _GEN_1082; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1084 = 4'h6 == _T_88695 ? shiftedStoreDataKnownPReg_6 : _GEN_1083; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1085 = 4'h7 == _T_88695 ? shiftedStoreDataKnownPReg_7 : _GEN_1084; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1086 = 4'h8 == _T_88695 ? shiftedStoreDataKnownPReg_8 : _GEN_1085; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1087 = 4'h9 == _T_88695 ? shiftedStoreDataKnownPReg_9 : _GEN_1086; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1088 = 4'ha == _T_88695 ? shiftedStoreDataKnownPReg_10 : _GEN_1087; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1089 = 4'hb == _T_88695 ? shiftedStoreDataKnownPReg_11 : _GEN_1088; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1090 = 4'hc == _T_88695 ? shiftedStoreDataKnownPReg_12 : _GEN_1089; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1091 = 4'hd == _T_88695 ? shiftedStoreDataKnownPReg_13 : _GEN_1090; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1092 = 4'he == _T_88695 ? shiftedStoreDataKnownPReg_14 : _GEN_1091; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1093 = 4'hf == _T_88695 ? shiftedStoreDataKnownPReg_15 : _GEN_1092; // @[AxiLoadQueue.scala 194:31:@35430.6]
  assign _GEN_1095 = 4'h1 == _T_88695 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1096 = 4'h2 == _T_88695 ? shiftedStoreDataQPreg_2 : _GEN_1095; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1097 = 4'h3 == _T_88695 ? shiftedStoreDataQPreg_3 : _GEN_1096; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1098 = 4'h4 == _T_88695 ? shiftedStoreDataQPreg_4 : _GEN_1097; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1099 = 4'h5 == _T_88695 ? shiftedStoreDataQPreg_5 : _GEN_1098; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1100 = 4'h6 == _T_88695 ? shiftedStoreDataQPreg_6 : _GEN_1099; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1101 = 4'h7 == _T_88695 ? shiftedStoreDataQPreg_7 : _GEN_1100; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1102 = 4'h8 == _T_88695 ? shiftedStoreDataQPreg_8 : _GEN_1101; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1103 = 4'h9 == _T_88695 ? shiftedStoreDataQPreg_9 : _GEN_1102; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1104 = 4'ha == _T_88695 ? shiftedStoreDataQPreg_10 : _GEN_1103; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1105 = 4'hb == _T_88695 ? shiftedStoreDataQPreg_11 : _GEN_1104; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1106 = 4'hc == _T_88695 ? shiftedStoreDataQPreg_12 : _GEN_1105; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1107 = 4'hd == _T_88695 ? shiftedStoreDataQPreg_13 : _GEN_1106; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1108 = 4'he == _T_88695 ? shiftedStoreDataQPreg_14 : _GEN_1107; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign _GEN_1109 = 4'hf == _T_88695 ? shiftedStoreDataQPreg_15 : _GEN_1108; // @[AxiLoadQueue.scala 195:31:@35431.6]
  assign lastConflict_3_0 = _T_88712 ? _GEN_1062 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_1 = _T_88712 ? _GEN_1063 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_2 = _T_88712 ? _GEN_1064 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_3 = _T_88712 ? _GEN_1065 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_4 = _T_88712 ? _GEN_1066 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_5 = _T_88712 ? _GEN_1067 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_6 = _T_88712 ? _GEN_1068 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_7 = _T_88712 ? _GEN_1069 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_8 = _T_88712 ? _GEN_1070 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_9 = _T_88712 ? _GEN_1071 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_10 = _T_88712 ? _GEN_1072 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_11 = _T_88712 ? _GEN_1073 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_12 = _T_88712 ? _GEN_1074 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_13 = _T_88712 ? _GEN_1075 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_14 = _T_88712 ? _GEN_1076 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign lastConflict_3_15 = _T_88712 ? _GEN_1077 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign canBypass_3 = _T_88712 ? _GEN_1093 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign bypassVal_3 = _T_88712 ? _GEN_1109 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35428.4]
  assign _T_88818 = conflictPReg_4_2 ? 2'h2 : {{1'd0}, conflictPReg_4_1}; // @[AxiLoadQueue.scala 191:60:@35485.4]
  assign _T_88819 = conflictPReg_4_3 ? 2'h3 : _T_88818; // @[AxiLoadQueue.scala 191:60:@35486.4]
  assign _T_88820 = conflictPReg_4_4 ? 3'h4 : {{1'd0}, _T_88819}; // @[AxiLoadQueue.scala 191:60:@35487.4]
  assign _T_88821 = conflictPReg_4_5 ? 3'h5 : _T_88820; // @[AxiLoadQueue.scala 191:60:@35488.4]
  assign _T_88822 = conflictPReg_4_6 ? 3'h6 : _T_88821; // @[AxiLoadQueue.scala 191:60:@35489.4]
  assign _T_88823 = conflictPReg_4_7 ? 3'h7 : _T_88822; // @[AxiLoadQueue.scala 191:60:@35490.4]
  assign _T_88824 = conflictPReg_4_8 ? 4'h8 : {{1'd0}, _T_88823}; // @[AxiLoadQueue.scala 191:60:@35491.4]
  assign _T_88825 = conflictPReg_4_9 ? 4'h9 : _T_88824; // @[AxiLoadQueue.scala 191:60:@35492.4]
  assign _T_88826 = conflictPReg_4_10 ? 4'ha : _T_88825; // @[AxiLoadQueue.scala 191:60:@35493.4]
  assign _T_88827 = conflictPReg_4_11 ? 4'hb : _T_88826; // @[AxiLoadQueue.scala 191:60:@35494.4]
  assign _T_88828 = conflictPReg_4_12 ? 4'hc : _T_88827; // @[AxiLoadQueue.scala 191:60:@35495.4]
  assign _T_88829 = conflictPReg_4_13 ? 4'hd : _T_88828; // @[AxiLoadQueue.scala 191:60:@35496.4]
  assign _T_88830 = conflictPReg_4_14 ? 4'he : _T_88829; // @[AxiLoadQueue.scala 191:60:@35497.4]
  assign _T_88831 = conflictPReg_4_15 ? 4'hf : _T_88830; // @[AxiLoadQueue.scala 191:60:@35498.4]
  assign _T_88834 = conflictPReg_4_0 | conflictPReg_4_1; // @[AxiLoadQueue.scala 192:43:@35500.4]
  assign _T_88835 = _T_88834 | conflictPReg_4_2; // @[AxiLoadQueue.scala 192:43:@35501.4]
  assign _T_88836 = _T_88835 | conflictPReg_4_3; // @[AxiLoadQueue.scala 192:43:@35502.4]
  assign _T_88837 = _T_88836 | conflictPReg_4_4; // @[AxiLoadQueue.scala 192:43:@35503.4]
  assign _T_88838 = _T_88837 | conflictPReg_4_5; // @[AxiLoadQueue.scala 192:43:@35504.4]
  assign _T_88839 = _T_88838 | conflictPReg_4_6; // @[AxiLoadQueue.scala 192:43:@35505.4]
  assign _T_88840 = _T_88839 | conflictPReg_4_7; // @[AxiLoadQueue.scala 192:43:@35506.4]
  assign _T_88841 = _T_88840 | conflictPReg_4_8; // @[AxiLoadQueue.scala 192:43:@35507.4]
  assign _T_88842 = _T_88841 | conflictPReg_4_9; // @[AxiLoadQueue.scala 192:43:@35508.4]
  assign _T_88843 = _T_88842 | conflictPReg_4_10; // @[AxiLoadQueue.scala 192:43:@35509.4]
  assign _T_88844 = _T_88843 | conflictPReg_4_11; // @[AxiLoadQueue.scala 192:43:@35510.4]
  assign _T_88845 = _T_88844 | conflictPReg_4_12; // @[AxiLoadQueue.scala 192:43:@35511.4]
  assign _T_88846 = _T_88845 | conflictPReg_4_13; // @[AxiLoadQueue.scala 192:43:@35512.4]
  assign _T_88847 = _T_88846 | conflictPReg_4_14; // @[AxiLoadQueue.scala 192:43:@35513.4]
  assign _T_88848 = _T_88847 | conflictPReg_4_15; // @[AxiLoadQueue.scala 192:43:@35514.4]
  assign _GEN_1128 = 4'h0 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1129 = 4'h1 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1130 = 4'h2 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1131 = 4'h3 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1132 = 4'h4 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1133 = 4'h5 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1134 = 4'h6 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1135 = 4'h7 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1136 = 4'h8 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1137 = 4'h9 == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1138 = 4'ha == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1139 = 4'hb == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1140 = 4'hc == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1141 = 4'hd == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1142 = 4'he == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1143 = 4'hf == _T_88831; // @[AxiLoadQueue.scala 193:43:@35516.6]
  assign _GEN_1145 = 4'h1 == _T_88831 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1146 = 4'h2 == _T_88831 ? shiftedStoreDataKnownPReg_2 : _GEN_1145; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1147 = 4'h3 == _T_88831 ? shiftedStoreDataKnownPReg_3 : _GEN_1146; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1148 = 4'h4 == _T_88831 ? shiftedStoreDataKnownPReg_4 : _GEN_1147; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1149 = 4'h5 == _T_88831 ? shiftedStoreDataKnownPReg_5 : _GEN_1148; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1150 = 4'h6 == _T_88831 ? shiftedStoreDataKnownPReg_6 : _GEN_1149; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1151 = 4'h7 == _T_88831 ? shiftedStoreDataKnownPReg_7 : _GEN_1150; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1152 = 4'h8 == _T_88831 ? shiftedStoreDataKnownPReg_8 : _GEN_1151; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1153 = 4'h9 == _T_88831 ? shiftedStoreDataKnownPReg_9 : _GEN_1152; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1154 = 4'ha == _T_88831 ? shiftedStoreDataKnownPReg_10 : _GEN_1153; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1155 = 4'hb == _T_88831 ? shiftedStoreDataKnownPReg_11 : _GEN_1154; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1156 = 4'hc == _T_88831 ? shiftedStoreDataKnownPReg_12 : _GEN_1155; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1157 = 4'hd == _T_88831 ? shiftedStoreDataKnownPReg_13 : _GEN_1156; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1158 = 4'he == _T_88831 ? shiftedStoreDataKnownPReg_14 : _GEN_1157; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1159 = 4'hf == _T_88831 ? shiftedStoreDataKnownPReg_15 : _GEN_1158; // @[AxiLoadQueue.scala 194:31:@35517.6]
  assign _GEN_1161 = 4'h1 == _T_88831 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1162 = 4'h2 == _T_88831 ? shiftedStoreDataQPreg_2 : _GEN_1161; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1163 = 4'h3 == _T_88831 ? shiftedStoreDataQPreg_3 : _GEN_1162; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1164 = 4'h4 == _T_88831 ? shiftedStoreDataQPreg_4 : _GEN_1163; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1165 = 4'h5 == _T_88831 ? shiftedStoreDataQPreg_5 : _GEN_1164; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1166 = 4'h6 == _T_88831 ? shiftedStoreDataQPreg_6 : _GEN_1165; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1167 = 4'h7 == _T_88831 ? shiftedStoreDataQPreg_7 : _GEN_1166; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1168 = 4'h8 == _T_88831 ? shiftedStoreDataQPreg_8 : _GEN_1167; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1169 = 4'h9 == _T_88831 ? shiftedStoreDataQPreg_9 : _GEN_1168; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1170 = 4'ha == _T_88831 ? shiftedStoreDataQPreg_10 : _GEN_1169; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1171 = 4'hb == _T_88831 ? shiftedStoreDataQPreg_11 : _GEN_1170; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1172 = 4'hc == _T_88831 ? shiftedStoreDataQPreg_12 : _GEN_1171; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1173 = 4'hd == _T_88831 ? shiftedStoreDataQPreg_13 : _GEN_1172; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1174 = 4'he == _T_88831 ? shiftedStoreDataQPreg_14 : _GEN_1173; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign _GEN_1175 = 4'hf == _T_88831 ? shiftedStoreDataQPreg_15 : _GEN_1174; // @[AxiLoadQueue.scala 195:31:@35518.6]
  assign lastConflict_4_0 = _T_88848 ? _GEN_1128 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_1 = _T_88848 ? _GEN_1129 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_2 = _T_88848 ? _GEN_1130 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_3 = _T_88848 ? _GEN_1131 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_4 = _T_88848 ? _GEN_1132 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_5 = _T_88848 ? _GEN_1133 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_6 = _T_88848 ? _GEN_1134 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_7 = _T_88848 ? _GEN_1135 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_8 = _T_88848 ? _GEN_1136 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_9 = _T_88848 ? _GEN_1137 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_10 = _T_88848 ? _GEN_1138 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_11 = _T_88848 ? _GEN_1139 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_12 = _T_88848 ? _GEN_1140 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_13 = _T_88848 ? _GEN_1141 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_14 = _T_88848 ? _GEN_1142 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign lastConflict_4_15 = _T_88848 ? _GEN_1143 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign canBypass_4 = _T_88848 ? _GEN_1159 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign bypassVal_4 = _T_88848 ? _GEN_1175 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35515.4]
  assign _T_88954 = conflictPReg_5_2 ? 2'h2 : {{1'd0}, conflictPReg_5_1}; // @[AxiLoadQueue.scala 191:60:@35572.4]
  assign _T_88955 = conflictPReg_5_3 ? 2'h3 : _T_88954; // @[AxiLoadQueue.scala 191:60:@35573.4]
  assign _T_88956 = conflictPReg_5_4 ? 3'h4 : {{1'd0}, _T_88955}; // @[AxiLoadQueue.scala 191:60:@35574.4]
  assign _T_88957 = conflictPReg_5_5 ? 3'h5 : _T_88956; // @[AxiLoadQueue.scala 191:60:@35575.4]
  assign _T_88958 = conflictPReg_5_6 ? 3'h6 : _T_88957; // @[AxiLoadQueue.scala 191:60:@35576.4]
  assign _T_88959 = conflictPReg_5_7 ? 3'h7 : _T_88958; // @[AxiLoadQueue.scala 191:60:@35577.4]
  assign _T_88960 = conflictPReg_5_8 ? 4'h8 : {{1'd0}, _T_88959}; // @[AxiLoadQueue.scala 191:60:@35578.4]
  assign _T_88961 = conflictPReg_5_9 ? 4'h9 : _T_88960; // @[AxiLoadQueue.scala 191:60:@35579.4]
  assign _T_88962 = conflictPReg_5_10 ? 4'ha : _T_88961; // @[AxiLoadQueue.scala 191:60:@35580.4]
  assign _T_88963 = conflictPReg_5_11 ? 4'hb : _T_88962; // @[AxiLoadQueue.scala 191:60:@35581.4]
  assign _T_88964 = conflictPReg_5_12 ? 4'hc : _T_88963; // @[AxiLoadQueue.scala 191:60:@35582.4]
  assign _T_88965 = conflictPReg_5_13 ? 4'hd : _T_88964; // @[AxiLoadQueue.scala 191:60:@35583.4]
  assign _T_88966 = conflictPReg_5_14 ? 4'he : _T_88965; // @[AxiLoadQueue.scala 191:60:@35584.4]
  assign _T_88967 = conflictPReg_5_15 ? 4'hf : _T_88966; // @[AxiLoadQueue.scala 191:60:@35585.4]
  assign _T_88970 = conflictPReg_5_0 | conflictPReg_5_1; // @[AxiLoadQueue.scala 192:43:@35587.4]
  assign _T_88971 = _T_88970 | conflictPReg_5_2; // @[AxiLoadQueue.scala 192:43:@35588.4]
  assign _T_88972 = _T_88971 | conflictPReg_5_3; // @[AxiLoadQueue.scala 192:43:@35589.4]
  assign _T_88973 = _T_88972 | conflictPReg_5_4; // @[AxiLoadQueue.scala 192:43:@35590.4]
  assign _T_88974 = _T_88973 | conflictPReg_5_5; // @[AxiLoadQueue.scala 192:43:@35591.4]
  assign _T_88975 = _T_88974 | conflictPReg_5_6; // @[AxiLoadQueue.scala 192:43:@35592.4]
  assign _T_88976 = _T_88975 | conflictPReg_5_7; // @[AxiLoadQueue.scala 192:43:@35593.4]
  assign _T_88977 = _T_88976 | conflictPReg_5_8; // @[AxiLoadQueue.scala 192:43:@35594.4]
  assign _T_88978 = _T_88977 | conflictPReg_5_9; // @[AxiLoadQueue.scala 192:43:@35595.4]
  assign _T_88979 = _T_88978 | conflictPReg_5_10; // @[AxiLoadQueue.scala 192:43:@35596.4]
  assign _T_88980 = _T_88979 | conflictPReg_5_11; // @[AxiLoadQueue.scala 192:43:@35597.4]
  assign _T_88981 = _T_88980 | conflictPReg_5_12; // @[AxiLoadQueue.scala 192:43:@35598.4]
  assign _T_88982 = _T_88981 | conflictPReg_5_13; // @[AxiLoadQueue.scala 192:43:@35599.4]
  assign _T_88983 = _T_88982 | conflictPReg_5_14; // @[AxiLoadQueue.scala 192:43:@35600.4]
  assign _T_88984 = _T_88983 | conflictPReg_5_15; // @[AxiLoadQueue.scala 192:43:@35601.4]
  assign _GEN_1194 = 4'h0 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1195 = 4'h1 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1196 = 4'h2 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1197 = 4'h3 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1198 = 4'h4 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1199 = 4'h5 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1200 = 4'h6 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1201 = 4'h7 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1202 = 4'h8 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1203 = 4'h9 == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1204 = 4'ha == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1205 = 4'hb == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1206 = 4'hc == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1207 = 4'hd == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1208 = 4'he == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1209 = 4'hf == _T_88967; // @[AxiLoadQueue.scala 193:43:@35603.6]
  assign _GEN_1211 = 4'h1 == _T_88967 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1212 = 4'h2 == _T_88967 ? shiftedStoreDataKnownPReg_2 : _GEN_1211; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1213 = 4'h3 == _T_88967 ? shiftedStoreDataKnownPReg_3 : _GEN_1212; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1214 = 4'h4 == _T_88967 ? shiftedStoreDataKnownPReg_4 : _GEN_1213; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1215 = 4'h5 == _T_88967 ? shiftedStoreDataKnownPReg_5 : _GEN_1214; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1216 = 4'h6 == _T_88967 ? shiftedStoreDataKnownPReg_6 : _GEN_1215; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1217 = 4'h7 == _T_88967 ? shiftedStoreDataKnownPReg_7 : _GEN_1216; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1218 = 4'h8 == _T_88967 ? shiftedStoreDataKnownPReg_8 : _GEN_1217; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1219 = 4'h9 == _T_88967 ? shiftedStoreDataKnownPReg_9 : _GEN_1218; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1220 = 4'ha == _T_88967 ? shiftedStoreDataKnownPReg_10 : _GEN_1219; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1221 = 4'hb == _T_88967 ? shiftedStoreDataKnownPReg_11 : _GEN_1220; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1222 = 4'hc == _T_88967 ? shiftedStoreDataKnownPReg_12 : _GEN_1221; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1223 = 4'hd == _T_88967 ? shiftedStoreDataKnownPReg_13 : _GEN_1222; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1224 = 4'he == _T_88967 ? shiftedStoreDataKnownPReg_14 : _GEN_1223; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1225 = 4'hf == _T_88967 ? shiftedStoreDataKnownPReg_15 : _GEN_1224; // @[AxiLoadQueue.scala 194:31:@35604.6]
  assign _GEN_1227 = 4'h1 == _T_88967 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1228 = 4'h2 == _T_88967 ? shiftedStoreDataQPreg_2 : _GEN_1227; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1229 = 4'h3 == _T_88967 ? shiftedStoreDataQPreg_3 : _GEN_1228; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1230 = 4'h4 == _T_88967 ? shiftedStoreDataQPreg_4 : _GEN_1229; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1231 = 4'h5 == _T_88967 ? shiftedStoreDataQPreg_5 : _GEN_1230; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1232 = 4'h6 == _T_88967 ? shiftedStoreDataQPreg_6 : _GEN_1231; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1233 = 4'h7 == _T_88967 ? shiftedStoreDataQPreg_7 : _GEN_1232; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1234 = 4'h8 == _T_88967 ? shiftedStoreDataQPreg_8 : _GEN_1233; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1235 = 4'h9 == _T_88967 ? shiftedStoreDataQPreg_9 : _GEN_1234; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1236 = 4'ha == _T_88967 ? shiftedStoreDataQPreg_10 : _GEN_1235; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1237 = 4'hb == _T_88967 ? shiftedStoreDataQPreg_11 : _GEN_1236; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1238 = 4'hc == _T_88967 ? shiftedStoreDataQPreg_12 : _GEN_1237; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1239 = 4'hd == _T_88967 ? shiftedStoreDataQPreg_13 : _GEN_1238; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1240 = 4'he == _T_88967 ? shiftedStoreDataQPreg_14 : _GEN_1239; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign _GEN_1241 = 4'hf == _T_88967 ? shiftedStoreDataQPreg_15 : _GEN_1240; // @[AxiLoadQueue.scala 195:31:@35605.6]
  assign lastConflict_5_0 = _T_88984 ? _GEN_1194 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_1 = _T_88984 ? _GEN_1195 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_2 = _T_88984 ? _GEN_1196 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_3 = _T_88984 ? _GEN_1197 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_4 = _T_88984 ? _GEN_1198 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_5 = _T_88984 ? _GEN_1199 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_6 = _T_88984 ? _GEN_1200 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_7 = _T_88984 ? _GEN_1201 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_8 = _T_88984 ? _GEN_1202 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_9 = _T_88984 ? _GEN_1203 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_10 = _T_88984 ? _GEN_1204 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_11 = _T_88984 ? _GEN_1205 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_12 = _T_88984 ? _GEN_1206 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_13 = _T_88984 ? _GEN_1207 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_14 = _T_88984 ? _GEN_1208 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign lastConflict_5_15 = _T_88984 ? _GEN_1209 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign canBypass_5 = _T_88984 ? _GEN_1225 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign bypassVal_5 = _T_88984 ? _GEN_1241 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35602.4]
  assign _T_89090 = conflictPReg_6_2 ? 2'h2 : {{1'd0}, conflictPReg_6_1}; // @[AxiLoadQueue.scala 191:60:@35659.4]
  assign _T_89091 = conflictPReg_6_3 ? 2'h3 : _T_89090; // @[AxiLoadQueue.scala 191:60:@35660.4]
  assign _T_89092 = conflictPReg_6_4 ? 3'h4 : {{1'd0}, _T_89091}; // @[AxiLoadQueue.scala 191:60:@35661.4]
  assign _T_89093 = conflictPReg_6_5 ? 3'h5 : _T_89092; // @[AxiLoadQueue.scala 191:60:@35662.4]
  assign _T_89094 = conflictPReg_6_6 ? 3'h6 : _T_89093; // @[AxiLoadQueue.scala 191:60:@35663.4]
  assign _T_89095 = conflictPReg_6_7 ? 3'h7 : _T_89094; // @[AxiLoadQueue.scala 191:60:@35664.4]
  assign _T_89096 = conflictPReg_6_8 ? 4'h8 : {{1'd0}, _T_89095}; // @[AxiLoadQueue.scala 191:60:@35665.4]
  assign _T_89097 = conflictPReg_6_9 ? 4'h9 : _T_89096; // @[AxiLoadQueue.scala 191:60:@35666.4]
  assign _T_89098 = conflictPReg_6_10 ? 4'ha : _T_89097; // @[AxiLoadQueue.scala 191:60:@35667.4]
  assign _T_89099 = conflictPReg_6_11 ? 4'hb : _T_89098; // @[AxiLoadQueue.scala 191:60:@35668.4]
  assign _T_89100 = conflictPReg_6_12 ? 4'hc : _T_89099; // @[AxiLoadQueue.scala 191:60:@35669.4]
  assign _T_89101 = conflictPReg_6_13 ? 4'hd : _T_89100; // @[AxiLoadQueue.scala 191:60:@35670.4]
  assign _T_89102 = conflictPReg_6_14 ? 4'he : _T_89101; // @[AxiLoadQueue.scala 191:60:@35671.4]
  assign _T_89103 = conflictPReg_6_15 ? 4'hf : _T_89102; // @[AxiLoadQueue.scala 191:60:@35672.4]
  assign _T_89106 = conflictPReg_6_0 | conflictPReg_6_1; // @[AxiLoadQueue.scala 192:43:@35674.4]
  assign _T_89107 = _T_89106 | conflictPReg_6_2; // @[AxiLoadQueue.scala 192:43:@35675.4]
  assign _T_89108 = _T_89107 | conflictPReg_6_3; // @[AxiLoadQueue.scala 192:43:@35676.4]
  assign _T_89109 = _T_89108 | conflictPReg_6_4; // @[AxiLoadQueue.scala 192:43:@35677.4]
  assign _T_89110 = _T_89109 | conflictPReg_6_5; // @[AxiLoadQueue.scala 192:43:@35678.4]
  assign _T_89111 = _T_89110 | conflictPReg_6_6; // @[AxiLoadQueue.scala 192:43:@35679.4]
  assign _T_89112 = _T_89111 | conflictPReg_6_7; // @[AxiLoadQueue.scala 192:43:@35680.4]
  assign _T_89113 = _T_89112 | conflictPReg_6_8; // @[AxiLoadQueue.scala 192:43:@35681.4]
  assign _T_89114 = _T_89113 | conflictPReg_6_9; // @[AxiLoadQueue.scala 192:43:@35682.4]
  assign _T_89115 = _T_89114 | conflictPReg_6_10; // @[AxiLoadQueue.scala 192:43:@35683.4]
  assign _T_89116 = _T_89115 | conflictPReg_6_11; // @[AxiLoadQueue.scala 192:43:@35684.4]
  assign _T_89117 = _T_89116 | conflictPReg_6_12; // @[AxiLoadQueue.scala 192:43:@35685.4]
  assign _T_89118 = _T_89117 | conflictPReg_6_13; // @[AxiLoadQueue.scala 192:43:@35686.4]
  assign _T_89119 = _T_89118 | conflictPReg_6_14; // @[AxiLoadQueue.scala 192:43:@35687.4]
  assign _T_89120 = _T_89119 | conflictPReg_6_15; // @[AxiLoadQueue.scala 192:43:@35688.4]
  assign _GEN_1260 = 4'h0 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1261 = 4'h1 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1262 = 4'h2 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1263 = 4'h3 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1264 = 4'h4 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1265 = 4'h5 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1266 = 4'h6 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1267 = 4'h7 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1268 = 4'h8 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1269 = 4'h9 == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1270 = 4'ha == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1271 = 4'hb == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1272 = 4'hc == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1273 = 4'hd == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1274 = 4'he == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1275 = 4'hf == _T_89103; // @[AxiLoadQueue.scala 193:43:@35690.6]
  assign _GEN_1277 = 4'h1 == _T_89103 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1278 = 4'h2 == _T_89103 ? shiftedStoreDataKnownPReg_2 : _GEN_1277; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1279 = 4'h3 == _T_89103 ? shiftedStoreDataKnownPReg_3 : _GEN_1278; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1280 = 4'h4 == _T_89103 ? shiftedStoreDataKnownPReg_4 : _GEN_1279; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1281 = 4'h5 == _T_89103 ? shiftedStoreDataKnownPReg_5 : _GEN_1280; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1282 = 4'h6 == _T_89103 ? shiftedStoreDataKnownPReg_6 : _GEN_1281; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1283 = 4'h7 == _T_89103 ? shiftedStoreDataKnownPReg_7 : _GEN_1282; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1284 = 4'h8 == _T_89103 ? shiftedStoreDataKnownPReg_8 : _GEN_1283; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1285 = 4'h9 == _T_89103 ? shiftedStoreDataKnownPReg_9 : _GEN_1284; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1286 = 4'ha == _T_89103 ? shiftedStoreDataKnownPReg_10 : _GEN_1285; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1287 = 4'hb == _T_89103 ? shiftedStoreDataKnownPReg_11 : _GEN_1286; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1288 = 4'hc == _T_89103 ? shiftedStoreDataKnownPReg_12 : _GEN_1287; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1289 = 4'hd == _T_89103 ? shiftedStoreDataKnownPReg_13 : _GEN_1288; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1290 = 4'he == _T_89103 ? shiftedStoreDataKnownPReg_14 : _GEN_1289; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1291 = 4'hf == _T_89103 ? shiftedStoreDataKnownPReg_15 : _GEN_1290; // @[AxiLoadQueue.scala 194:31:@35691.6]
  assign _GEN_1293 = 4'h1 == _T_89103 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1294 = 4'h2 == _T_89103 ? shiftedStoreDataQPreg_2 : _GEN_1293; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1295 = 4'h3 == _T_89103 ? shiftedStoreDataQPreg_3 : _GEN_1294; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1296 = 4'h4 == _T_89103 ? shiftedStoreDataQPreg_4 : _GEN_1295; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1297 = 4'h5 == _T_89103 ? shiftedStoreDataQPreg_5 : _GEN_1296; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1298 = 4'h6 == _T_89103 ? shiftedStoreDataQPreg_6 : _GEN_1297; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1299 = 4'h7 == _T_89103 ? shiftedStoreDataQPreg_7 : _GEN_1298; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1300 = 4'h8 == _T_89103 ? shiftedStoreDataQPreg_8 : _GEN_1299; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1301 = 4'h9 == _T_89103 ? shiftedStoreDataQPreg_9 : _GEN_1300; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1302 = 4'ha == _T_89103 ? shiftedStoreDataQPreg_10 : _GEN_1301; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1303 = 4'hb == _T_89103 ? shiftedStoreDataQPreg_11 : _GEN_1302; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1304 = 4'hc == _T_89103 ? shiftedStoreDataQPreg_12 : _GEN_1303; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1305 = 4'hd == _T_89103 ? shiftedStoreDataQPreg_13 : _GEN_1304; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1306 = 4'he == _T_89103 ? shiftedStoreDataQPreg_14 : _GEN_1305; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign _GEN_1307 = 4'hf == _T_89103 ? shiftedStoreDataQPreg_15 : _GEN_1306; // @[AxiLoadQueue.scala 195:31:@35692.6]
  assign lastConflict_6_0 = _T_89120 ? _GEN_1260 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_1 = _T_89120 ? _GEN_1261 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_2 = _T_89120 ? _GEN_1262 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_3 = _T_89120 ? _GEN_1263 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_4 = _T_89120 ? _GEN_1264 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_5 = _T_89120 ? _GEN_1265 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_6 = _T_89120 ? _GEN_1266 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_7 = _T_89120 ? _GEN_1267 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_8 = _T_89120 ? _GEN_1268 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_9 = _T_89120 ? _GEN_1269 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_10 = _T_89120 ? _GEN_1270 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_11 = _T_89120 ? _GEN_1271 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_12 = _T_89120 ? _GEN_1272 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_13 = _T_89120 ? _GEN_1273 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_14 = _T_89120 ? _GEN_1274 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign lastConflict_6_15 = _T_89120 ? _GEN_1275 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign canBypass_6 = _T_89120 ? _GEN_1291 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign bypassVal_6 = _T_89120 ? _GEN_1307 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35689.4]
  assign _T_89226 = conflictPReg_7_2 ? 2'h2 : {{1'd0}, conflictPReg_7_1}; // @[AxiLoadQueue.scala 191:60:@35746.4]
  assign _T_89227 = conflictPReg_7_3 ? 2'h3 : _T_89226; // @[AxiLoadQueue.scala 191:60:@35747.4]
  assign _T_89228 = conflictPReg_7_4 ? 3'h4 : {{1'd0}, _T_89227}; // @[AxiLoadQueue.scala 191:60:@35748.4]
  assign _T_89229 = conflictPReg_7_5 ? 3'h5 : _T_89228; // @[AxiLoadQueue.scala 191:60:@35749.4]
  assign _T_89230 = conflictPReg_7_6 ? 3'h6 : _T_89229; // @[AxiLoadQueue.scala 191:60:@35750.4]
  assign _T_89231 = conflictPReg_7_7 ? 3'h7 : _T_89230; // @[AxiLoadQueue.scala 191:60:@35751.4]
  assign _T_89232 = conflictPReg_7_8 ? 4'h8 : {{1'd0}, _T_89231}; // @[AxiLoadQueue.scala 191:60:@35752.4]
  assign _T_89233 = conflictPReg_7_9 ? 4'h9 : _T_89232; // @[AxiLoadQueue.scala 191:60:@35753.4]
  assign _T_89234 = conflictPReg_7_10 ? 4'ha : _T_89233; // @[AxiLoadQueue.scala 191:60:@35754.4]
  assign _T_89235 = conflictPReg_7_11 ? 4'hb : _T_89234; // @[AxiLoadQueue.scala 191:60:@35755.4]
  assign _T_89236 = conflictPReg_7_12 ? 4'hc : _T_89235; // @[AxiLoadQueue.scala 191:60:@35756.4]
  assign _T_89237 = conflictPReg_7_13 ? 4'hd : _T_89236; // @[AxiLoadQueue.scala 191:60:@35757.4]
  assign _T_89238 = conflictPReg_7_14 ? 4'he : _T_89237; // @[AxiLoadQueue.scala 191:60:@35758.4]
  assign _T_89239 = conflictPReg_7_15 ? 4'hf : _T_89238; // @[AxiLoadQueue.scala 191:60:@35759.4]
  assign _T_89242 = conflictPReg_7_0 | conflictPReg_7_1; // @[AxiLoadQueue.scala 192:43:@35761.4]
  assign _T_89243 = _T_89242 | conflictPReg_7_2; // @[AxiLoadQueue.scala 192:43:@35762.4]
  assign _T_89244 = _T_89243 | conflictPReg_7_3; // @[AxiLoadQueue.scala 192:43:@35763.4]
  assign _T_89245 = _T_89244 | conflictPReg_7_4; // @[AxiLoadQueue.scala 192:43:@35764.4]
  assign _T_89246 = _T_89245 | conflictPReg_7_5; // @[AxiLoadQueue.scala 192:43:@35765.4]
  assign _T_89247 = _T_89246 | conflictPReg_7_6; // @[AxiLoadQueue.scala 192:43:@35766.4]
  assign _T_89248 = _T_89247 | conflictPReg_7_7; // @[AxiLoadQueue.scala 192:43:@35767.4]
  assign _T_89249 = _T_89248 | conflictPReg_7_8; // @[AxiLoadQueue.scala 192:43:@35768.4]
  assign _T_89250 = _T_89249 | conflictPReg_7_9; // @[AxiLoadQueue.scala 192:43:@35769.4]
  assign _T_89251 = _T_89250 | conflictPReg_7_10; // @[AxiLoadQueue.scala 192:43:@35770.4]
  assign _T_89252 = _T_89251 | conflictPReg_7_11; // @[AxiLoadQueue.scala 192:43:@35771.4]
  assign _T_89253 = _T_89252 | conflictPReg_7_12; // @[AxiLoadQueue.scala 192:43:@35772.4]
  assign _T_89254 = _T_89253 | conflictPReg_7_13; // @[AxiLoadQueue.scala 192:43:@35773.4]
  assign _T_89255 = _T_89254 | conflictPReg_7_14; // @[AxiLoadQueue.scala 192:43:@35774.4]
  assign _T_89256 = _T_89255 | conflictPReg_7_15; // @[AxiLoadQueue.scala 192:43:@35775.4]
  assign _GEN_1326 = 4'h0 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1327 = 4'h1 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1328 = 4'h2 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1329 = 4'h3 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1330 = 4'h4 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1331 = 4'h5 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1332 = 4'h6 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1333 = 4'h7 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1334 = 4'h8 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1335 = 4'h9 == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1336 = 4'ha == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1337 = 4'hb == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1338 = 4'hc == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1339 = 4'hd == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1340 = 4'he == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1341 = 4'hf == _T_89239; // @[AxiLoadQueue.scala 193:43:@35777.6]
  assign _GEN_1343 = 4'h1 == _T_89239 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1344 = 4'h2 == _T_89239 ? shiftedStoreDataKnownPReg_2 : _GEN_1343; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1345 = 4'h3 == _T_89239 ? shiftedStoreDataKnownPReg_3 : _GEN_1344; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1346 = 4'h4 == _T_89239 ? shiftedStoreDataKnownPReg_4 : _GEN_1345; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1347 = 4'h5 == _T_89239 ? shiftedStoreDataKnownPReg_5 : _GEN_1346; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1348 = 4'h6 == _T_89239 ? shiftedStoreDataKnownPReg_6 : _GEN_1347; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1349 = 4'h7 == _T_89239 ? shiftedStoreDataKnownPReg_7 : _GEN_1348; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1350 = 4'h8 == _T_89239 ? shiftedStoreDataKnownPReg_8 : _GEN_1349; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1351 = 4'h9 == _T_89239 ? shiftedStoreDataKnownPReg_9 : _GEN_1350; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1352 = 4'ha == _T_89239 ? shiftedStoreDataKnownPReg_10 : _GEN_1351; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1353 = 4'hb == _T_89239 ? shiftedStoreDataKnownPReg_11 : _GEN_1352; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1354 = 4'hc == _T_89239 ? shiftedStoreDataKnownPReg_12 : _GEN_1353; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1355 = 4'hd == _T_89239 ? shiftedStoreDataKnownPReg_13 : _GEN_1354; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1356 = 4'he == _T_89239 ? shiftedStoreDataKnownPReg_14 : _GEN_1355; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1357 = 4'hf == _T_89239 ? shiftedStoreDataKnownPReg_15 : _GEN_1356; // @[AxiLoadQueue.scala 194:31:@35778.6]
  assign _GEN_1359 = 4'h1 == _T_89239 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1360 = 4'h2 == _T_89239 ? shiftedStoreDataQPreg_2 : _GEN_1359; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1361 = 4'h3 == _T_89239 ? shiftedStoreDataQPreg_3 : _GEN_1360; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1362 = 4'h4 == _T_89239 ? shiftedStoreDataQPreg_4 : _GEN_1361; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1363 = 4'h5 == _T_89239 ? shiftedStoreDataQPreg_5 : _GEN_1362; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1364 = 4'h6 == _T_89239 ? shiftedStoreDataQPreg_6 : _GEN_1363; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1365 = 4'h7 == _T_89239 ? shiftedStoreDataQPreg_7 : _GEN_1364; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1366 = 4'h8 == _T_89239 ? shiftedStoreDataQPreg_8 : _GEN_1365; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1367 = 4'h9 == _T_89239 ? shiftedStoreDataQPreg_9 : _GEN_1366; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1368 = 4'ha == _T_89239 ? shiftedStoreDataQPreg_10 : _GEN_1367; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1369 = 4'hb == _T_89239 ? shiftedStoreDataQPreg_11 : _GEN_1368; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1370 = 4'hc == _T_89239 ? shiftedStoreDataQPreg_12 : _GEN_1369; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1371 = 4'hd == _T_89239 ? shiftedStoreDataQPreg_13 : _GEN_1370; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1372 = 4'he == _T_89239 ? shiftedStoreDataQPreg_14 : _GEN_1371; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign _GEN_1373 = 4'hf == _T_89239 ? shiftedStoreDataQPreg_15 : _GEN_1372; // @[AxiLoadQueue.scala 195:31:@35779.6]
  assign lastConflict_7_0 = _T_89256 ? _GEN_1326 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_1 = _T_89256 ? _GEN_1327 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_2 = _T_89256 ? _GEN_1328 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_3 = _T_89256 ? _GEN_1329 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_4 = _T_89256 ? _GEN_1330 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_5 = _T_89256 ? _GEN_1331 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_6 = _T_89256 ? _GEN_1332 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_7 = _T_89256 ? _GEN_1333 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_8 = _T_89256 ? _GEN_1334 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_9 = _T_89256 ? _GEN_1335 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_10 = _T_89256 ? _GEN_1336 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_11 = _T_89256 ? _GEN_1337 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_12 = _T_89256 ? _GEN_1338 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_13 = _T_89256 ? _GEN_1339 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_14 = _T_89256 ? _GEN_1340 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign lastConflict_7_15 = _T_89256 ? _GEN_1341 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign canBypass_7 = _T_89256 ? _GEN_1357 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign bypassVal_7 = _T_89256 ? _GEN_1373 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35776.4]
  assign _T_89362 = conflictPReg_8_2 ? 2'h2 : {{1'd0}, conflictPReg_8_1}; // @[AxiLoadQueue.scala 191:60:@35833.4]
  assign _T_89363 = conflictPReg_8_3 ? 2'h3 : _T_89362; // @[AxiLoadQueue.scala 191:60:@35834.4]
  assign _T_89364 = conflictPReg_8_4 ? 3'h4 : {{1'd0}, _T_89363}; // @[AxiLoadQueue.scala 191:60:@35835.4]
  assign _T_89365 = conflictPReg_8_5 ? 3'h5 : _T_89364; // @[AxiLoadQueue.scala 191:60:@35836.4]
  assign _T_89366 = conflictPReg_8_6 ? 3'h6 : _T_89365; // @[AxiLoadQueue.scala 191:60:@35837.4]
  assign _T_89367 = conflictPReg_8_7 ? 3'h7 : _T_89366; // @[AxiLoadQueue.scala 191:60:@35838.4]
  assign _T_89368 = conflictPReg_8_8 ? 4'h8 : {{1'd0}, _T_89367}; // @[AxiLoadQueue.scala 191:60:@35839.4]
  assign _T_89369 = conflictPReg_8_9 ? 4'h9 : _T_89368; // @[AxiLoadQueue.scala 191:60:@35840.4]
  assign _T_89370 = conflictPReg_8_10 ? 4'ha : _T_89369; // @[AxiLoadQueue.scala 191:60:@35841.4]
  assign _T_89371 = conflictPReg_8_11 ? 4'hb : _T_89370; // @[AxiLoadQueue.scala 191:60:@35842.4]
  assign _T_89372 = conflictPReg_8_12 ? 4'hc : _T_89371; // @[AxiLoadQueue.scala 191:60:@35843.4]
  assign _T_89373 = conflictPReg_8_13 ? 4'hd : _T_89372; // @[AxiLoadQueue.scala 191:60:@35844.4]
  assign _T_89374 = conflictPReg_8_14 ? 4'he : _T_89373; // @[AxiLoadQueue.scala 191:60:@35845.4]
  assign _T_89375 = conflictPReg_8_15 ? 4'hf : _T_89374; // @[AxiLoadQueue.scala 191:60:@35846.4]
  assign _T_89378 = conflictPReg_8_0 | conflictPReg_8_1; // @[AxiLoadQueue.scala 192:43:@35848.4]
  assign _T_89379 = _T_89378 | conflictPReg_8_2; // @[AxiLoadQueue.scala 192:43:@35849.4]
  assign _T_89380 = _T_89379 | conflictPReg_8_3; // @[AxiLoadQueue.scala 192:43:@35850.4]
  assign _T_89381 = _T_89380 | conflictPReg_8_4; // @[AxiLoadQueue.scala 192:43:@35851.4]
  assign _T_89382 = _T_89381 | conflictPReg_8_5; // @[AxiLoadQueue.scala 192:43:@35852.4]
  assign _T_89383 = _T_89382 | conflictPReg_8_6; // @[AxiLoadQueue.scala 192:43:@35853.4]
  assign _T_89384 = _T_89383 | conflictPReg_8_7; // @[AxiLoadQueue.scala 192:43:@35854.4]
  assign _T_89385 = _T_89384 | conflictPReg_8_8; // @[AxiLoadQueue.scala 192:43:@35855.4]
  assign _T_89386 = _T_89385 | conflictPReg_8_9; // @[AxiLoadQueue.scala 192:43:@35856.4]
  assign _T_89387 = _T_89386 | conflictPReg_8_10; // @[AxiLoadQueue.scala 192:43:@35857.4]
  assign _T_89388 = _T_89387 | conflictPReg_8_11; // @[AxiLoadQueue.scala 192:43:@35858.4]
  assign _T_89389 = _T_89388 | conflictPReg_8_12; // @[AxiLoadQueue.scala 192:43:@35859.4]
  assign _T_89390 = _T_89389 | conflictPReg_8_13; // @[AxiLoadQueue.scala 192:43:@35860.4]
  assign _T_89391 = _T_89390 | conflictPReg_8_14; // @[AxiLoadQueue.scala 192:43:@35861.4]
  assign _T_89392 = _T_89391 | conflictPReg_8_15; // @[AxiLoadQueue.scala 192:43:@35862.4]
  assign _GEN_1392 = 4'h0 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1393 = 4'h1 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1394 = 4'h2 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1395 = 4'h3 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1396 = 4'h4 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1397 = 4'h5 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1398 = 4'h6 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1399 = 4'h7 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1400 = 4'h8 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1401 = 4'h9 == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1402 = 4'ha == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1403 = 4'hb == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1404 = 4'hc == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1405 = 4'hd == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1406 = 4'he == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1407 = 4'hf == _T_89375; // @[AxiLoadQueue.scala 193:43:@35864.6]
  assign _GEN_1409 = 4'h1 == _T_89375 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1410 = 4'h2 == _T_89375 ? shiftedStoreDataKnownPReg_2 : _GEN_1409; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1411 = 4'h3 == _T_89375 ? shiftedStoreDataKnownPReg_3 : _GEN_1410; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1412 = 4'h4 == _T_89375 ? shiftedStoreDataKnownPReg_4 : _GEN_1411; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1413 = 4'h5 == _T_89375 ? shiftedStoreDataKnownPReg_5 : _GEN_1412; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1414 = 4'h6 == _T_89375 ? shiftedStoreDataKnownPReg_6 : _GEN_1413; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1415 = 4'h7 == _T_89375 ? shiftedStoreDataKnownPReg_7 : _GEN_1414; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1416 = 4'h8 == _T_89375 ? shiftedStoreDataKnownPReg_8 : _GEN_1415; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1417 = 4'h9 == _T_89375 ? shiftedStoreDataKnownPReg_9 : _GEN_1416; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1418 = 4'ha == _T_89375 ? shiftedStoreDataKnownPReg_10 : _GEN_1417; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1419 = 4'hb == _T_89375 ? shiftedStoreDataKnownPReg_11 : _GEN_1418; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1420 = 4'hc == _T_89375 ? shiftedStoreDataKnownPReg_12 : _GEN_1419; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1421 = 4'hd == _T_89375 ? shiftedStoreDataKnownPReg_13 : _GEN_1420; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1422 = 4'he == _T_89375 ? shiftedStoreDataKnownPReg_14 : _GEN_1421; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1423 = 4'hf == _T_89375 ? shiftedStoreDataKnownPReg_15 : _GEN_1422; // @[AxiLoadQueue.scala 194:31:@35865.6]
  assign _GEN_1425 = 4'h1 == _T_89375 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1426 = 4'h2 == _T_89375 ? shiftedStoreDataQPreg_2 : _GEN_1425; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1427 = 4'h3 == _T_89375 ? shiftedStoreDataQPreg_3 : _GEN_1426; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1428 = 4'h4 == _T_89375 ? shiftedStoreDataQPreg_4 : _GEN_1427; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1429 = 4'h5 == _T_89375 ? shiftedStoreDataQPreg_5 : _GEN_1428; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1430 = 4'h6 == _T_89375 ? shiftedStoreDataQPreg_6 : _GEN_1429; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1431 = 4'h7 == _T_89375 ? shiftedStoreDataQPreg_7 : _GEN_1430; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1432 = 4'h8 == _T_89375 ? shiftedStoreDataQPreg_8 : _GEN_1431; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1433 = 4'h9 == _T_89375 ? shiftedStoreDataQPreg_9 : _GEN_1432; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1434 = 4'ha == _T_89375 ? shiftedStoreDataQPreg_10 : _GEN_1433; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1435 = 4'hb == _T_89375 ? shiftedStoreDataQPreg_11 : _GEN_1434; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1436 = 4'hc == _T_89375 ? shiftedStoreDataQPreg_12 : _GEN_1435; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1437 = 4'hd == _T_89375 ? shiftedStoreDataQPreg_13 : _GEN_1436; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1438 = 4'he == _T_89375 ? shiftedStoreDataQPreg_14 : _GEN_1437; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign _GEN_1439 = 4'hf == _T_89375 ? shiftedStoreDataQPreg_15 : _GEN_1438; // @[AxiLoadQueue.scala 195:31:@35866.6]
  assign lastConflict_8_0 = _T_89392 ? _GEN_1392 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_1 = _T_89392 ? _GEN_1393 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_2 = _T_89392 ? _GEN_1394 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_3 = _T_89392 ? _GEN_1395 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_4 = _T_89392 ? _GEN_1396 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_5 = _T_89392 ? _GEN_1397 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_6 = _T_89392 ? _GEN_1398 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_7 = _T_89392 ? _GEN_1399 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_8 = _T_89392 ? _GEN_1400 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_9 = _T_89392 ? _GEN_1401 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_10 = _T_89392 ? _GEN_1402 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_11 = _T_89392 ? _GEN_1403 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_12 = _T_89392 ? _GEN_1404 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_13 = _T_89392 ? _GEN_1405 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_14 = _T_89392 ? _GEN_1406 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign lastConflict_8_15 = _T_89392 ? _GEN_1407 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign canBypass_8 = _T_89392 ? _GEN_1423 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign bypassVal_8 = _T_89392 ? _GEN_1439 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35863.4]
  assign _T_89498 = conflictPReg_9_2 ? 2'h2 : {{1'd0}, conflictPReg_9_1}; // @[AxiLoadQueue.scala 191:60:@35920.4]
  assign _T_89499 = conflictPReg_9_3 ? 2'h3 : _T_89498; // @[AxiLoadQueue.scala 191:60:@35921.4]
  assign _T_89500 = conflictPReg_9_4 ? 3'h4 : {{1'd0}, _T_89499}; // @[AxiLoadQueue.scala 191:60:@35922.4]
  assign _T_89501 = conflictPReg_9_5 ? 3'h5 : _T_89500; // @[AxiLoadQueue.scala 191:60:@35923.4]
  assign _T_89502 = conflictPReg_9_6 ? 3'h6 : _T_89501; // @[AxiLoadQueue.scala 191:60:@35924.4]
  assign _T_89503 = conflictPReg_9_7 ? 3'h7 : _T_89502; // @[AxiLoadQueue.scala 191:60:@35925.4]
  assign _T_89504 = conflictPReg_9_8 ? 4'h8 : {{1'd0}, _T_89503}; // @[AxiLoadQueue.scala 191:60:@35926.4]
  assign _T_89505 = conflictPReg_9_9 ? 4'h9 : _T_89504; // @[AxiLoadQueue.scala 191:60:@35927.4]
  assign _T_89506 = conflictPReg_9_10 ? 4'ha : _T_89505; // @[AxiLoadQueue.scala 191:60:@35928.4]
  assign _T_89507 = conflictPReg_9_11 ? 4'hb : _T_89506; // @[AxiLoadQueue.scala 191:60:@35929.4]
  assign _T_89508 = conflictPReg_9_12 ? 4'hc : _T_89507; // @[AxiLoadQueue.scala 191:60:@35930.4]
  assign _T_89509 = conflictPReg_9_13 ? 4'hd : _T_89508; // @[AxiLoadQueue.scala 191:60:@35931.4]
  assign _T_89510 = conflictPReg_9_14 ? 4'he : _T_89509; // @[AxiLoadQueue.scala 191:60:@35932.4]
  assign _T_89511 = conflictPReg_9_15 ? 4'hf : _T_89510; // @[AxiLoadQueue.scala 191:60:@35933.4]
  assign _T_89514 = conflictPReg_9_0 | conflictPReg_9_1; // @[AxiLoadQueue.scala 192:43:@35935.4]
  assign _T_89515 = _T_89514 | conflictPReg_9_2; // @[AxiLoadQueue.scala 192:43:@35936.4]
  assign _T_89516 = _T_89515 | conflictPReg_9_3; // @[AxiLoadQueue.scala 192:43:@35937.4]
  assign _T_89517 = _T_89516 | conflictPReg_9_4; // @[AxiLoadQueue.scala 192:43:@35938.4]
  assign _T_89518 = _T_89517 | conflictPReg_9_5; // @[AxiLoadQueue.scala 192:43:@35939.4]
  assign _T_89519 = _T_89518 | conflictPReg_9_6; // @[AxiLoadQueue.scala 192:43:@35940.4]
  assign _T_89520 = _T_89519 | conflictPReg_9_7; // @[AxiLoadQueue.scala 192:43:@35941.4]
  assign _T_89521 = _T_89520 | conflictPReg_9_8; // @[AxiLoadQueue.scala 192:43:@35942.4]
  assign _T_89522 = _T_89521 | conflictPReg_9_9; // @[AxiLoadQueue.scala 192:43:@35943.4]
  assign _T_89523 = _T_89522 | conflictPReg_9_10; // @[AxiLoadQueue.scala 192:43:@35944.4]
  assign _T_89524 = _T_89523 | conflictPReg_9_11; // @[AxiLoadQueue.scala 192:43:@35945.4]
  assign _T_89525 = _T_89524 | conflictPReg_9_12; // @[AxiLoadQueue.scala 192:43:@35946.4]
  assign _T_89526 = _T_89525 | conflictPReg_9_13; // @[AxiLoadQueue.scala 192:43:@35947.4]
  assign _T_89527 = _T_89526 | conflictPReg_9_14; // @[AxiLoadQueue.scala 192:43:@35948.4]
  assign _T_89528 = _T_89527 | conflictPReg_9_15; // @[AxiLoadQueue.scala 192:43:@35949.4]
  assign _GEN_1458 = 4'h0 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1459 = 4'h1 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1460 = 4'h2 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1461 = 4'h3 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1462 = 4'h4 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1463 = 4'h5 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1464 = 4'h6 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1465 = 4'h7 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1466 = 4'h8 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1467 = 4'h9 == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1468 = 4'ha == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1469 = 4'hb == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1470 = 4'hc == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1471 = 4'hd == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1472 = 4'he == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1473 = 4'hf == _T_89511; // @[AxiLoadQueue.scala 193:43:@35951.6]
  assign _GEN_1475 = 4'h1 == _T_89511 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1476 = 4'h2 == _T_89511 ? shiftedStoreDataKnownPReg_2 : _GEN_1475; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1477 = 4'h3 == _T_89511 ? shiftedStoreDataKnownPReg_3 : _GEN_1476; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1478 = 4'h4 == _T_89511 ? shiftedStoreDataKnownPReg_4 : _GEN_1477; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1479 = 4'h5 == _T_89511 ? shiftedStoreDataKnownPReg_5 : _GEN_1478; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1480 = 4'h6 == _T_89511 ? shiftedStoreDataKnownPReg_6 : _GEN_1479; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1481 = 4'h7 == _T_89511 ? shiftedStoreDataKnownPReg_7 : _GEN_1480; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1482 = 4'h8 == _T_89511 ? shiftedStoreDataKnownPReg_8 : _GEN_1481; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1483 = 4'h9 == _T_89511 ? shiftedStoreDataKnownPReg_9 : _GEN_1482; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1484 = 4'ha == _T_89511 ? shiftedStoreDataKnownPReg_10 : _GEN_1483; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1485 = 4'hb == _T_89511 ? shiftedStoreDataKnownPReg_11 : _GEN_1484; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1486 = 4'hc == _T_89511 ? shiftedStoreDataKnownPReg_12 : _GEN_1485; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1487 = 4'hd == _T_89511 ? shiftedStoreDataKnownPReg_13 : _GEN_1486; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1488 = 4'he == _T_89511 ? shiftedStoreDataKnownPReg_14 : _GEN_1487; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1489 = 4'hf == _T_89511 ? shiftedStoreDataKnownPReg_15 : _GEN_1488; // @[AxiLoadQueue.scala 194:31:@35952.6]
  assign _GEN_1491 = 4'h1 == _T_89511 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1492 = 4'h2 == _T_89511 ? shiftedStoreDataQPreg_2 : _GEN_1491; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1493 = 4'h3 == _T_89511 ? shiftedStoreDataQPreg_3 : _GEN_1492; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1494 = 4'h4 == _T_89511 ? shiftedStoreDataQPreg_4 : _GEN_1493; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1495 = 4'h5 == _T_89511 ? shiftedStoreDataQPreg_5 : _GEN_1494; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1496 = 4'h6 == _T_89511 ? shiftedStoreDataQPreg_6 : _GEN_1495; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1497 = 4'h7 == _T_89511 ? shiftedStoreDataQPreg_7 : _GEN_1496; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1498 = 4'h8 == _T_89511 ? shiftedStoreDataQPreg_8 : _GEN_1497; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1499 = 4'h9 == _T_89511 ? shiftedStoreDataQPreg_9 : _GEN_1498; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1500 = 4'ha == _T_89511 ? shiftedStoreDataQPreg_10 : _GEN_1499; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1501 = 4'hb == _T_89511 ? shiftedStoreDataQPreg_11 : _GEN_1500; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1502 = 4'hc == _T_89511 ? shiftedStoreDataQPreg_12 : _GEN_1501; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1503 = 4'hd == _T_89511 ? shiftedStoreDataQPreg_13 : _GEN_1502; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1504 = 4'he == _T_89511 ? shiftedStoreDataQPreg_14 : _GEN_1503; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign _GEN_1505 = 4'hf == _T_89511 ? shiftedStoreDataQPreg_15 : _GEN_1504; // @[AxiLoadQueue.scala 195:31:@35953.6]
  assign lastConflict_9_0 = _T_89528 ? _GEN_1458 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_1 = _T_89528 ? _GEN_1459 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_2 = _T_89528 ? _GEN_1460 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_3 = _T_89528 ? _GEN_1461 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_4 = _T_89528 ? _GEN_1462 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_5 = _T_89528 ? _GEN_1463 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_6 = _T_89528 ? _GEN_1464 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_7 = _T_89528 ? _GEN_1465 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_8 = _T_89528 ? _GEN_1466 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_9 = _T_89528 ? _GEN_1467 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_10 = _T_89528 ? _GEN_1468 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_11 = _T_89528 ? _GEN_1469 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_12 = _T_89528 ? _GEN_1470 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_13 = _T_89528 ? _GEN_1471 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_14 = _T_89528 ? _GEN_1472 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign lastConflict_9_15 = _T_89528 ? _GEN_1473 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign canBypass_9 = _T_89528 ? _GEN_1489 : 1'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign bypassVal_9 = _T_89528 ? _GEN_1505 : 32'h0; // @[AxiLoadQueue.scala 192:53:@35950.4]
  assign _T_89634 = conflictPReg_10_2 ? 2'h2 : {{1'd0}, conflictPReg_10_1}; // @[AxiLoadQueue.scala 191:60:@36007.4]
  assign _T_89635 = conflictPReg_10_3 ? 2'h3 : _T_89634; // @[AxiLoadQueue.scala 191:60:@36008.4]
  assign _T_89636 = conflictPReg_10_4 ? 3'h4 : {{1'd0}, _T_89635}; // @[AxiLoadQueue.scala 191:60:@36009.4]
  assign _T_89637 = conflictPReg_10_5 ? 3'h5 : _T_89636; // @[AxiLoadQueue.scala 191:60:@36010.4]
  assign _T_89638 = conflictPReg_10_6 ? 3'h6 : _T_89637; // @[AxiLoadQueue.scala 191:60:@36011.4]
  assign _T_89639 = conflictPReg_10_7 ? 3'h7 : _T_89638; // @[AxiLoadQueue.scala 191:60:@36012.4]
  assign _T_89640 = conflictPReg_10_8 ? 4'h8 : {{1'd0}, _T_89639}; // @[AxiLoadQueue.scala 191:60:@36013.4]
  assign _T_89641 = conflictPReg_10_9 ? 4'h9 : _T_89640; // @[AxiLoadQueue.scala 191:60:@36014.4]
  assign _T_89642 = conflictPReg_10_10 ? 4'ha : _T_89641; // @[AxiLoadQueue.scala 191:60:@36015.4]
  assign _T_89643 = conflictPReg_10_11 ? 4'hb : _T_89642; // @[AxiLoadQueue.scala 191:60:@36016.4]
  assign _T_89644 = conflictPReg_10_12 ? 4'hc : _T_89643; // @[AxiLoadQueue.scala 191:60:@36017.4]
  assign _T_89645 = conflictPReg_10_13 ? 4'hd : _T_89644; // @[AxiLoadQueue.scala 191:60:@36018.4]
  assign _T_89646 = conflictPReg_10_14 ? 4'he : _T_89645; // @[AxiLoadQueue.scala 191:60:@36019.4]
  assign _T_89647 = conflictPReg_10_15 ? 4'hf : _T_89646; // @[AxiLoadQueue.scala 191:60:@36020.4]
  assign _T_89650 = conflictPReg_10_0 | conflictPReg_10_1; // @[AxiLoadQueue.scala 192:43:@36022.4]
  assign _T_89651 = _T_89650 | conflictPReg_10_2; // @[AxiLoadQueue.scala 192:43:@36023.4]
  assign _T_89652 = _T_89651 | conflictPReg_10_3; // @[AxiLoadQueue.scala 192:43:@36024.4]
  assign _T_89653 = _T_89652 | conflictPReg_10_4; // @[AxiLoadQueue.scala 192:43:@36025.4]
  assign _T_89654 = _T_89653 | conflictPReg_10_5; // @[AxiLoadQueue.scala 192:43:@36026.4]
  assign _T_89655 = _T_89654 | conflictPReg_10_6; // @[AxiLoadQueue.scala 192:43:@36027.4]
  assign _T_89656 = _T_89655 | conflictPReg_10_7; // @[AxiLoadQueue.scala 192:43:@36028.4]
  assign _T_89657 = _T_89656 | conflictPReg_10_8; // @[AxiLoadQueue.scala 192:43:@36029.4]
  assign _T_89658 = _T_89657 | conflictPReg_10_9; // @[AxiLoadQueue.scala 192:43:@36030.4]
  assign _T_89659 = _T_89658 | conflictPReg_10_10; // @[AxiLoadQueue.scala 192:43:@36031.4]
  assign _T_89660 = _T_89659 | conflictPReg_10_11; // @[AxiLoadQueue.scala 192:43:@36032.4]
  assign _T_89661 = _T_89660 | conflictPReg_10_12; // @[AxiLoadQueue.scala 192:43:@36033.4]
  assign _T_89662 = _T_89661 | conflictPReg_10_13; // @[AxiLoadQueue.scala 192:43:@36034.4]
  assign _T_89663 = _T_89662 | conflictPReg_10_14; // @[AxiLoadQueue.scala 192:43:@36035.4]
  assign _T_89664 = _T_89663 | conflictPReg_10_15; // @[AxiLoadQueue.scala 192:43:@36036.4]
  assign _GEN_1524 = 4'h0 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1525 = 4'h1 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1526 = 4'h2 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1527 = 4'h3 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1528 = 4'h4 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1529 = 4'h5 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1530 = 4'h6 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1531 = 4'h7 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1532 = 4'h8 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1533 = 4'h9 == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1534 = 4'ha == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1535 = 4'hb == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1536 = 4'hc == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1537 = 4'hd == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1538 = 4'he == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1539 = 4'hf == _T_89647; // @[AxiLoadQueue.scala 193:43:@36038.6]
  assign _GEN_1541 = 4'h1 == _T_89647 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1542 = 4'h2 == _T_89647 ? shiftedStoreDataKnownPReg_2 : _GEN_1541; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1543 = 4'h3 == _T_89647 ? shiftedStoreDataKnownPReg_3 : _GEN_1542; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1544 = 4'h4 == _T_89647 ? shiftedStoreDataKnownPReg_4 : _GEN_1543; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1545 = 4'h5 == _T_89647 ? shiftedStoreDataKnownPReg_5 : _GEN_1544; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1546 = 4'h6 == _T_89647 ? shiftedStoreDataKnownPReg_6 : _GEN_1545; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1547 = 4'h7 == _T_89647 ? shiftedStoreDataKnownPReg_7 : _GEN_1546; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1548 = 4'h8 == _T_89647 ? shiftedStoreDataKnownPReg_8 : _GEN_1547; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1549 = 4'h9 == _T_89647 ? shiftedStoreDataKnownPReg_9 : _GEN_1548; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1550 = 4'ha == _T_89647 ? shiftedStoreDataKnownPReg_10 : _GEN_1549; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1551 = 4'hb == _T_89647 ? shiftedStoreDataKnownPReg_11 : _GEN_1550; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1552 = 4'hc == _T_89647 ? shiftedStoreDataKnownPReg_12 : _GEN_1551; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1553 = 4'hd == _T_89647 ? shiftedStoreDataKnownPReg_13 : _GEN_1552; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1554 = 4'he == _T_89647 ? shiftedStoreDataKnownPReg_14 : _GEN_1553; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1555 = 4'hf == _T_89647 ? shiftedStoreDataKnownPReg_15 : _GEN_1554; // @[AxiLoadQueue.scala 194:31:@36039.6]
  assign _GEN_1557 = 4'h1 == _T_89647 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1558 = 4'h2 == _T_89647 ? shiftedStoreDataQPreg_2 : _GEN_1557; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1559 = 4'h3 == _T_89647 ? shiftedStoreDataQPreg_3 : _GEN_1558; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1560 = 4'h4 == _T_89647 ? shiftedStoreDataQPreg_4 : _GEN_1559; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1561 = 4'h5 == _T_89647 ? shiftedStoreDataQPreg_5 : _GEN_1560; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1562 = 4'h6 == _T_89647 ? shiftedStoreDataQPreg_6 : _GEN_1561; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1563 = 4'h7 == _T_89647 ? shiftedStoreDataQPreg_7 : _GEN_1562; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1564 = 4'h8 == _T_89647 ? shiftedStoreDataQPreg_8 : _GEN_1563; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1565 = 4'h9 == _T_89647 ? shiftedStoreDataQPreg_9 : _GEN_1564; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1566 = 4'ha == _T_89647 ? shiftedStoreDataQPreg_10 : _GEN_1565; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1567 = 4'hb == _T_89647 ? shiftedStoreDataQPreg_11 : _GEN_1566; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1568 = 4'hc == _T_89647 ? shiftedStoreDataQPreg_12 : _GEN_1567; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1569 = 4'hd == _T_89647 ? shiftedStoreDataQPreg_13 : _GEN_1568; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1570 = 4'he == _T_89647 ? shiftedStoreDataQPreg_14 : _GEN_1569; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign _GEN_1571 = 4'hf == _T_89647 ? shiftedStoreDataQPreg_15 : _GEN_1570; // @[AxiLoadQueue.scala 195:31:@36040.6]
  assign lastConflict_10_0 = _T_89664 ? _GEN_1524 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_1 = _T_89664 ? _GEN_1525 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_2 = _T_89664 ? _GEN_1526 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_3 = _T_89664 ? _GEN_1527 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_4 = _T_89664 ? _GEN_1528 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_5 = _T_89664 ? _GEN_1529 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_6 = _T_89664 ? _GEN_1530 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_7 = _T_89664 ? _GEN_1531 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_8 = _T_89664 ? _GEN_1532 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_9 = _T_89664 ? _GEN_1533 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_10 = _T_89664 ? _GEN_1534 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_11 = _T_89664 ? _GEN_1535 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_12 = _T_89664 ? _GEN_1536 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_13 = _T_89664 ? _GEN_1537 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_14 = _T_89664 ? _GEN_1538 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign lastConflict_10_15 = _T_89664 ? _GEN_1539 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign canBypass_10 = _T_89664 ? _GEN_1555 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign bypassVal_10 = _T_89664 ? _GEN_1571 : 32'h0; // @[AxiLoadQueue.scala 192:53:@36037.4]
  assign _T_89770 = conflictPReg_11_2 ? 2'h2 : {{1'd0}, conflictPReg_11_1}; // @[AxiLoadQueue.scala 191:60:@36094.4]
  assign _T_89771 = conflictPReg_11_3 ? 2'h3 : _T_89770; // @[AxiLoadQueue.scala 191:60:@36095.4]
  assign _T_89772 = conflictPReg_11_4 ? 3'h4 : {{1'd0}, _T_89771}; // @[AxiLoadQueue.scala 191:60:@36096.4]
  assign _T_89773 = conflictPReg_11_5 ? 3'h5 : _T_89772; // @[AxiLoadQueue.scala 191:60:@36097.4]
  assign _T_89774 = conflictPReg_11_6 ? 3'h6 : _T_89773; // @[AxiLoadQueue.scala 191:60:@36098.4]
  assign _T_89775 = conflictPReg_11_7 ? 3'h7 : _T_89774; // @[AxiLoadQueue.scala 191:60:@36099.4]
  assign _T_89776 = conflictPReg_11_8 ? 4'h8 : {{1'd0}, _T_89775}; // @[AxiLoadQueue.scala 191:60:@36100.4]
  assign _T_89777 = conflictPReg_11_9 ? 4'h9 : _T_89776; // @[AxiLoadQueue.scala 191:60:@36101.4]
  assign _T_89778 = conflictPReg_11_10 ? 4'ha : _T_89777; // @[AxiLoadQueue.scala 191:60:@36102.4]
  assign _T_89779 = conflictPReg_11_11 ? 4'hb : _T_89778; // @[AxiLoadQueue.scala 191:60:@36103.4]
  assign _T_89780 = conflictPReg_11_12 ? 4'hc : _T_89779; // @[AxiLoadQueue.scala 191:60:@36104.4]
  assign _T_89781 = conflictPReg_11_13 ? 4'hd : _T_89780; // @[AxiLoadQueue.scala 191:60:@36105.4]
  assign _T_89782 = conflictPReg_11_14 ? 4'he : _T_89781; // @[AxiLoadQueue.scala 191:60:@36106.4]
  assign _T_89783 = conflictPReg_11_15 ? 4'hf : _T_89782; // @[AxiLoadQueue.scala 191:60:@36107.4]
  assign _T_89786 = conflictPReg_11_0 | conflictPReg_11_1; // @[AxiLoadQueue.scala 192:43:@36109.4]
  assign _T_89787 = _T_89786 | conflictPReg_11_2; // @[AxiLoadQueue.scala 192:43:@36110.4]
  assign _T_89788 = _T_89787 | conflictPReg_11_3; // @[AxiLoadQueue.scala 192:43:@36111.4]
  assign _T_89789 = _T_89788 | conflictPReg_11_4; // @[AxiLoadQueue.scala 192:43:@36112.4]
  assign _T_89790 = _T_89789 | conflictPReg_11_5; // @[AxiLoadQueue.scala 192:43:@36113.4]
  assign _T_89791 = _T_89790 | conflictPReg_11_6; // @[AxiLoadQueue.scala 192:43:@36114.4]
  assign _T_89792 = _T_89791 | conflictPReg_11_7; // @[AxiLoadQueue.scala 192:43:@36115.4]
  assign _T_89793 = _T_89792 | conflictPReg_11_8; // @[AxiLoadQueue.scala 192:43:@36116.4]
  assign _T_89794 = _T_89793 | conflictPReg_11_9; // @[AxiLoadQueue.scala 192:43:@36117.4]
  assign _T_89795 = _T_89794 | conflictPReg_11_10; // @[AxiLoadQueue.scala 192:43:@36118.4]
  assign _T_89796 = _T_89795 | conflictPReg_11_11; // @[AxiLoadQueue.scala 192:43:@36119.4]
  assign _T_89797 = _T_89796 | conflictPReg_11_12; // @[AxiLoadQueue.scala 192:43:@36120.4]
  assign _T_89798 = _T_89797 | conflictPReg_11_13; // @[AxiLoadQueue.scala 192:43:@36121.4]
  assign _T_89799 = _T_89798 | conflictPReg_11_14; // @[AxiLoadQueue.scala 192:43:@36122.4]
  assign _T_89800 = _T_89799 | conflictPReg_11_15; // @[AxiLoadQueue.scala 192:43:@36123.4]
  assign _GEN_1590 = 4'h0 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1591 = 4'h1 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1592 = 4'h2 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1593 = 4'h3 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1594 = 4'h4 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1595 = 4'h5 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1596 = 4'h6 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1597 = 4'h7 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1598 = 4'h8 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1599 = 4'h9 == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1600 = 4'ha == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1601 = 4'hb == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1602 = 4'hc == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1603 = 4'hd == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1604 = 4'he == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1605 = 4'hf == _T_89783; // @[AxiLoadQueue.scala 193:43:@36125.6]
  assign _GEN_1607 = 4'h1 == _T_89783 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1608 = 4'h2 == _T_89783 ? shiftedStoreDataKnownPReg_2 : _GEN_1607; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1609 = 4'h3 == _T_89783 ? shiftedStoreDataKnownPReg_3 : _GEN_1608; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1610 = 4'h4 == _T_89783 ? shiftedStoreDataKnownPReg_4 : _GEN_1609; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1611 = 4'h5 == _T_89783 ? shiftedStoreDataKnownPReg_5 : _GEN_1610; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1612 = 4'h6 == _T_89783 ? shiftedStoreDataKnownPReg_6 : _GEN_1611; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1613 = 4'h7 == _T_89783 ? shiftedStoreDataKnownPReg_7 : _GEN_1612; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1614 = 4'h8 == _T_89783 ? shiftedStoreDataKnownPReg_8 : _GEN_1613; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1615 = 4'h9 == _T_89783 ? shiftedStoreDataKnownPReg_9 : _GEN_1614; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1616 = 4'ha == _T_89783 ? shiftedStoreDataKnownPReg_10 : _GEN_1615; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1617 = 4'hb == _T_89783 ? shiftedStoreDataKnownPReg_11 : _GEN_1616; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1618 = 4'hc == _T_89783 ? shiftedStoreDataKnownPReg_12 : _GEN_1617; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1619 = 4'hd == _T_89783 ? shiftedStoreDataKnownPReg_13 : _GEN_1618; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1620 = 4'he == _T_89783 ? shiftedStoreDataKnownPReg_14 : _GEN_1619; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1621 = 4'hf == _T_89783 ? shiftedStoreDataKnownPReg_15 : _GEN_1620; // @[AxiLoadQueue.scala 194:31:@36126.6]
  assign _GEN_1623 = 4'h1 == _T_89783 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1624 = 4'h2 == _T_89783 ? shiftedStoreDataQPreg_2 : _GEN_1623; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1625 = 4'h3 == _T_89783 ? shiftedStoreDataQPreg_3 : _GEN_1624; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1626 = 4'h4 == _T_89783 ? shiftedStoreDataQPreg_4 : _GEN_1625; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1627 = 4'h5 == _T_89783 ? shiftedStoreDataQPreg_5 : _GEN_1626; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1628 = 4'h6 == _T_89783 ? shiftedStoreDataQPreg_6 : _GEN_1627; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1629 = 4'h7 == _T_89783 ? shiftedStoreDataQPreg_7 : _GEN_1628; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1630 = 4'h8 == _T_89783 ? shiftedStoreDataQPreg_8 : _GEN_1629; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1631 = 4'h9 == _T_89783 ? shiftedStoreDataQPreg_9 : _GEN_1630; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1632 = 4'ha == _T_89783 ? shiftedStoreDataQPreg_10 : _GEN_1631; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1633 = 4'hb == _T_89783 ? shiftedStoreDataQPreg_11 : _GEN_1632; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1634 = 4'hc == _T_89783 ? shiftedStoreDataQPreg_12 : _GEN_1633; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1635 = 4'hd == _T_89783 ? shiftedStoreDataQPreg_13 : _GEN_1634; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1636 = 4'he == _T_89783 ? shiftedStoreDataQPreg_14 : _GEN_1635; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign _GEN_1637 = 4'hf == _T_89783 ? shiftedStoreDataQPreg_15 : _GEN_1636; // @[AxiLoadQueue.scala 195:31:@36127.6]
  assign lastConflict_11_0 = _T_89800 ? _GEN_1590 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_1 = _T_89800 ? _GEN_1591 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_2 = _T_89800 ? _GEN_1592 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_3 = _T_89800 ? _GEN_1593 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_4 = _T_89800 ? _GEN_1594 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_5 = _T_89800 ? _GEN_1595 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_6 = _T_89800 ? _GEN_1596 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_7 = _T_89800 ? _GEN_1597 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_8 = _T_89800 ? _GEN_1598 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_9 = _T_89800 ? _GEN_1599 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_10 = _T_89800 ? _GEN_1600 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_11 = _T_89800 ? _GEN_1601 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_12 = _T_89800 ? _GEN_1602 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_13 = _T_89800 ? _GEN_1603 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_14 = _T_89800 ? _GEN_1604 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign lastConflict_11_15 = _T_89800 ? _GEN_1605 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign canBypass_11 = _T_89800 ? _GEN_1621 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign bypassVal_11 = _T_89800 ? _GEN_1637 : 32'h0; // @[AxiLoadQueue.scala 192:53:@36124.4]
  assign _T_89906 = conflictPReg_12_2 ? 2'h2 : {{1'd0}, conflictPReg_12_1}; // @[AxiLoadQueue.scala 191:60:@36181.4]
  assign _T_89907 = conflictPReg_12_3 ? 2'h3 : _T_89906; // @[AxiLoadQueue.scala 191:60:@36182.4]
  assign _T_89908 = conflictPReg_12_4 ? 3'h4 : {{1'd0}, _T_89907}; // @[AxiLoadQueue.scala 191:60:@36183.4]
  assign _T_89909 = conflictPReg_12_5 ? 3'h5 : _T_89908; // @[AxiLoadQueue.scala 191:60:@36184.4]
  assign _T_89910 = conflictPReg_12_6 ? 3'h6 : _T_89909; // @[AxiLoadQueue.scala 191:60:@36185.4]
  assign _T_89911 = conflictPReg_12_7 ? 3'h7 : _T_89910; // @[AxiLoadQueue.scala 191:60:@36186.4]
  assign _T_89912 = conflictPReg_12_8 ? 4'h8 : {{1'd0}, _T_89911}; // @[AxiLoadQueue.scala 191:60:@36187.4]
  assign _T_89913 = conflictPReg_12_9 ? 4'h9 : _T_89912; // @[AxiLoadQueue.scala 191:60:@36188.4]
  assign _T_89914 = conflictPReg_12_10 ? 4'ha : _T_89913; // @[AxiLoadQueue.scala 191:60:@36189.4]
  assign _T_89915 = conflictPReg_12_11 ? 4'hb : _T_89914; // @[AxiLoadQueue.scala 191:60:@36190.4]
  assign _T_89916 = conflictPReg_12_12 ? 4'hc : _T_89915; // @[AxiLoadQueue.scala 191:60:@36191.4]
  assign _T_89917 = conflictPReg_12_13 ? 4'hd : _T_89916; // @[AxiLoadQueue.scala 191:60:@36192.4]
  assign _T_89918 = conflictPReg_12_14 ? 4'he : _T_89917; // @[AxiLoadQueue.scala 191:60:@36193.4]
  assign _T_89919 = conflictPReg_12_15 ? 4'hf : _T_89918; // @[AxiLoadQueue.scala 191:60:@36194.4]
  assign _T_89922 = conflictPReg_12_0 | conflictPReg_12_1; // @[AxiLoadQueue.scala 192:43:@36196.4]
  assign _T_89923 = _T_89922 | conflictPReg_12_2; // @[AxiLoadQueue.scala 192:43:@36197.4]
  assign _T_89924 = _T_89923 | conflictPReg_12_3; // @[AxiLoadQueue.scala 192:43:@36198.4]
  assign _T_89925 = _T_89924 | conflictPReg_12_4; // @[AxiLoadQueue.scala 192:43:@36199.4]
  assign _T_89926 = _T_89925 | conflictPReg_12_5; // @[AxiLoadQueue.scala 192:43:@36200.4]
  assign _T_89927 = _T_89926 | conflictPReg_12_6; // @[AxiLoadQueue.scala 192:43:@36201.4]
  assign _T_89928 = _T_89927 | conflictPReg_12_7; // @[AxiLoadQueue.scala 192:43:@36202.4]
  assign _T_89929 = _T_89928 | conflictPReg_12_8; // @[AxiLoadQueue.scala 192:43:@36203.4]
  assign _T_89930 = _T_89929 | conflictPReg_12_9; // @[AxiLoadQueue.scala 192:43:@36204.4]
  assign _T_89931 = _T_89930 | conflictPReg_12_10; // @[AxiLoadQueue.scala 192:43:@36205.4]
  assign _T_89932 = _T_89931 | conflictPReg_12_11; // @[AxiLoadQueue.scala 192:43:@36206.4]
  assign _T_89933 = _T_89932 | conflictPReg_12_12; // @[AxiLoadQueue.scala 192:43:@36207.4]
  assign _T_89934 = _T_89933 | conflictPReg_12_13; // @[AxiLoadQueue.scala 192:43:@36208.4]
  assign _T_89935 = _T_89934 | conflictPReg_12_14; // @[AxiLoadQueue.scala 192:43:@36209.4]
  assign _T_89936 = _T_89935 | conflictPReg_12_15; // @[AxiLoadQueue.scala 192:43:@36210.4]
  assign _GEN_1656 = 4'h0 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1657 = 4'h1 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1658 = 4'h2 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1659 = 4'h3 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1660 = 4'h4 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1661 = 4'h5 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1662 = 4'h6 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1663 = 4'h7 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1664 = 4'h8 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1665 = 4'h9 == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1666 = 4'ha == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1667 = 4'hb == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1668 = 4'hc == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1669 = 4'hd == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1670 = 4'he == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1671 = 4'hf == _T_89919; // @[AxiLoadQueue.scala 193:43:@36212.6]
  assign _GEN_1673 = 4'h1 == _T_89919 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1674 = 4'h2 == _T_89919 ? shiftedStoreDataKnownPReg_2 : _GEN_1673; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1675 = 4'h3 == _T_89919 ? shiftedStoreDataKnownPReg_3 : _GEN_1674; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1676 = 4'h4 == _T_89919 ? shiftedStoreDataKnownPReg_4 : _GEN_1675; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1677 = 4'h5 == _T_89919 ? shiftedStoreDataKnownPReg_5 : _GEN_1676; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1678 = 4'h6 == _T_89919 ? shiftedStoreDataKnownPReg_6 : _GEN_1677; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1679 = 4'h7 == _T_89919 ? shiftedStoreDataKnownPReg_7 : _GEN_1678; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1680 = 4'h8 == _T_89919 ? shiftedStoreDataKnownPReg_8 : _GEN_1679; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1681 = 4'h9 == _T_89919 ? shiftedStoreDataKnownPReg_9 : _GEN_1680; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1682 = 4'ha == _T_89919 ? shiftedStoreDataKnownPReg_10 : _GEN_1681; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1683 = 4'hb == _T_89919 ? shiftedStoreDataKnownPReg_11 : _GEN_1682; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1684 = 4'hc == _T_89919 ? shiftedStoreDataKnownPReg_12 : _GEN_1683; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1685 = 4'hd == _T_89919 ? shiftedStoreDataKnownPReg_13 : _GEN_1684; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1686 = 4'he == _T_89919 ? shiftedStoreDataKnownPReg_14 : _GEN_1685; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1687 = 4'hf == _T_89919 ? shiftedStoreDataKnownPReg_15 : _GEN_1686; // @[AxiLoadQueue.scala 194:31:@36213.6]
  assign _GEN_1689 = 4'h1 == _T_89919 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1690 = 4'h2 == _T_89919 ? shiftedStoreDataQPreg_2 : _GEN_1689; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1691 = 4'h3 == _T_89919 ? shiftedStoreDataQPreg_3 : _GEN_1690; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1692 = 4'h4 == _T_89919 ? shiftedStoreDataQPreg_4 : _GEN_1691; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1693 = 4'h5 == _T_89919 ? shiftedStoreDataQPreg_5 : _GEN_1692; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1694 = 4'h6 == _T_89919 ? shiftedStoreDataQPreg_6 : _GEN_1693; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1695 = 4'h7 == _T_89919 ? shiftedStoreDataQPreg_7 : _GEN_1694; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1696 = 4'h8 == _T_89919 ? shiftedStoreDataQPreg_8 : _GEN_1695; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1697 = 4'h9 == _T_89919 ? shiftedStoreDataQPreg_9 : _GEN_1696; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1698 = 4'ha == _T_89919 ? shiftedStoreDataQPreg_10 : _GEN_1697; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1699 = 4'hb == _T_89919 ? shiftedStoreDataQPreg_11 : _GEN_1698; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1700 = 4'hc == _T_89919 ? shiftedStoreDataQPreg_12 : _GEN_1699; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1701 = 4'hd == _T_89919 ? shiftedStoreDataQPreg_13 : _GEN_1700; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1702 = 4'he == _T_89919 ? shiftedStoreDataQPreg_14 : _GEN_1701; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign _GEN_1703 = 4'hf == _T_89919 ? shiftedStoreDataQPreg_15 : _GEN_1702; // @[AxiLoadQueue.scala 195:31:@36214.6]
  assign lastConflict_12_0 = _T_89936 ? _GEN_1656 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_1 = _T_89936 ? _GEN_1657 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_2 = _T_89936 ? _GEN_1658 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_3 = _T_89936 ? _GEN_1659 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_4 = _T_89936 ? _GEN_1660 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_5 = _T_89936 ? _GEN_1661 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_6 = _T_89936 ? _GEN_1662 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_7 = _T_89936 ? _GEN_1663 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_8 = _T_89936 ? _GEN_1664 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_9 = _T_89936 ? _GEN_1665 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_10 = _T_89936 ? _GEN_1666 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_11 = _T_89936 ? _GEN_1667 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_12 = _T_89936 ? _GEN_1668 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_13 = _T_89936 ? _GEN_1669 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_14 = _T_89936 ? _GEN_1670 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign lastConflict_12_15 = _T_89936 ? _GEN_1671 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign canBypass_12 = _T_89936 ? _GEN_1687 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign bypassVal_12 = _T_89936 ? _GEN_1703 : 32'h0; // @[AxiLoadQueue.scala 192:53:@36211.4]
  assign _T_90042 = conflictPReg_13_2 ? 2'h2 : {{1'd0}, conflictPReg_13_1}; // @[AxiLoadQueue.scala 191:60:@36268.4]
  assign _T_90043 = conflictPReg_13_3 ? 2'h3 : _T_90042; // @[AxiLoadQueue.scala 191:60:@36269.4]
  assign _T_90044 = conflictPReg_13_4 ? 3'h4 : {{1'd0}, _T_90043}; // @[AxiLoadQueue.scala 191:60:@36270.4]
  assign _T_90045 = conflictPReg_13_5 ? 3'h5 : _T_90044; // @[AxiLoadQueue.scala 191:60:@36271.4]
  assign _T_90046 = conflictPReg_13_6 ? 3'h6 : _T_90045; // @[AxiLoadQueue.scala 191:60:@36272.4]
  assign _T_90047 = conflictPReg_13_7 ? 3'h7 : _T_90046; // @[AxiLoadQueue.scala 191:60:@36273.4]
  assign _T_90048 = conflictPReg_13_8 ? 4'h8 : {{1'd0}, _T_90047}; // @[AxiLoadQueue.scala 191:60:@36274.4]
  assign _T_90049 = conflictPReg_13_9 ? 4'h9 : _T_90048; // @[AxiLoadQueue.scala 191:60:@36275.4]
  assign _T_90050 = conflictPReg_13_10 ? 4'ha : _T_90049; // @[AxiLoadQueue.scala 191:60:@36276.4]
  assign _T_90051 = conflictPReg_13_11 ? 4'hb : _T_90050; // @[AxiLoadQueue.scala 191:60:@36277.4]
  assign _T_90052 = conflictPReg_13_12 ? 4'hc : _T_90051; // @[AxiLoadQueue.scala 191:60:@36278.4]
  assign _T_90053 = conflictPReg_13_13 ? 4'hd : _T_90052; // @[AxiLoadQueue.scala 191:60:@36279.4]
  assign _T_90054 = conflictPReg_13_14 ? 4'he : _T_90053; // @[AxiLoadQueue.scala 191:60:@36280.4]
  assign _T_90055 = conflictPReg_13_15 ? 4'hf : _T_90054; // @[AxiLoadQueue.scala 191:60:@36281.4]
  assign _T_90058 = conflictPReg_13_0 | conflictPReg_13_1; // @[AxiLoadQueue.scala 192:43:@36283.4]
  assign _T_90059 = _T_90058 | conflictPReg_13_2; // @[AxiLoadQueue.scala 192:43:@36284.4]
  assign _T_90060 = _T_90059 | conflictPReg_13_3; // @[AxiLoadQueue.scala 192:43:@36285.4]
  assign _T_90061 = _T_90060 | conflictPReg_13_4; // @[AxiLoadQueue.scala 192:43:@36286.4]
  assign _T_90062 = _T_90061 | conflictPReg_13_5; // @[AxiLoadQueue.scala 192:43:@36287.4]
  assign _T_90063 = _T_90062 | conflictPReg_13_6; // @[AxiLoadQueue.scala 192:43:@36288.4]
  assign _T_90064 = _T_90063 | conflictPReg_13_7; // @[AxiLoadQueue.scala 192:43:@36289.4]
  assign _T_90065 = _T_90064 | conflictPReg_13_8; // @[AxiLoadQueue.scala 192:43:@36290.4]
  assign _T_90066 = _T_90065 | conflictPReg_13_9; // @[AxiLoadQueue.scala 192:43:@36291.4]
  assign _T_90067 = _T_90066 | conflictPReg_13_10; // @[AxiLoadQueue.scala 192:43:@36292.4]
  assign _T_90068 = _T_90067 | conflictPReg_13_11; // @[AxiLoadQueue.scala 192:43:@36293.4]
  assign _T_90069 = _T_90068 | conflictPReg_13_12; // @[AxiLoadQueue.scala 192:43:@36294.4]
  assign _T_90070 = _T_90069 | conflictPReg_13_13; // @[AxiLoadQueue.scala 192:43:@36295.4]
  assign _T_90071 = _T_90070 | conflictPReg_13_14; // @[AxiLoadQueue.scala 192:43:@36296.4]
  assign _T_90072 = _T_90071 | conflictPReg_13_15; // @[AxiLoadQueue.scala 192:43:@36297.4]
  assign _GEN_1722 = 4'h0 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1723 = 4'h1 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1724 = 4'h2 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1725 = 4'h3 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1726 = 4'h4 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1727 = 4'h5 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1728 = 4'h6 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1729 = 4'h7 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1730 = 4'h8 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1731 = 4'h9 == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1732 = 4'ha == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1733 = 4'hb == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1734 = 4'hc == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1735 = 4'hd == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1736 = 4'he == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1737 = 4'hf == _T_90055; // @[AxiLoadQueue.scala 193:43:@36299.6]
  assign _GEN_1739 = 4'h1 == _T_90055 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1740 = 4'h2 == _T_90055 ? shiftedStoreDataKnownPReg_2 : _GEN_1739; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1741 = 4'h3 == _T_90055 ? shiftedStoreDataKnownPReg_3 : _GEN_1740; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1742 = 4'h4 == _T_90055 ? shiftedStoreDataKnownPReg_4 : _GEN_1741; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1743 = 4'h5 == _T_90055 ? shiftedStoreDataKnownPReg_5 : _GEN_1742; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1744 = 4'h6 == _T_90055 ? shiftedStoreDataKnownPReg_6 : _GEN_1743; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1745 = 4'h7 == _T_90055 ? shiftedStoreDataKnownPReg_7 : _GEN_1744; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1746 = 4'h8 == _T_90055 ? shiftedStoreDataKnownPReg_8 : _GEN_1745; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1747 = 4'h9 == _T_90055 ? shiftedStoreDataKnownPReg_9 : _GEN_1746; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1748 = 4'ha == _T_90055 ? shiftedStoreDataKnownPReg_10 : _GEN_1747; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1749 = 4'hb == _T_90055 ? shiftedStoreDataKnownPReg_11 : _GEN_1748; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1750 = 4'hc == _T_90055 ? shiftedStoreDataKnownPReg_12 : _GEN_1749; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1751 = 4'hd == _T_90055 ? shiftedStoreDataKnownPReg_13 : _GEN_1750; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1752 = 4'he == _T_90055 ? shiftedStoreDataKnownPReg_14 : _GEN_1751; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1753 = 4'hf == _T_90055 ? shiftedStoreDataKnownPReg_15 : _GEN_1752; // @[AxiLoadQueue.scala 194:31:@36300.6]
  assign _GEN_1755 = 4'h1 == _T_90055 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1756 = 4'h2 == _T_90055 ? shiftedStoreDataQPreg_2 : _GEN_1755; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1757 = 4'h3 == _T_90055 ? shiftedStoreDataQPreg_3 : _GEN_1756; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1758 = 4'h4 == _T_90055 ? shiftedStoreDataQPreg_4 : _GEN_1757; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1759 = 4'h5 == _T_90055 ? shiftedStoreDataQPreg_5 : _GEN_1758; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1760 = 4'h6 == _T_90055 ? shiftedStoreDataQPreg_6 : _GEN_1759; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1761 = 4'h7 == _T_90055 ? shiftedStoreDataQPreg_7 : _GEN_1760; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1762 = 4'h8 == _T_90055 ? shiftedStoreDataQPreg_8 : _GEN_1761; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1763 = 4'h9 == _T_90055 ? shiftedStoreDataQPreg_9 : _GEN_1762; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1764 = 4'ha == _T_90055 ? shiftedStoreDataQPreg_10 : _GEN_1763; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1765 = 4'hb == _T_90055 ? shiftedStoreDataQPreg_11 : _GEN_1764; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1766 = 4'hc == _T_90055 ? shiftedStoreDataQPreg_12 : _GEN_1765; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1767 = 4'hd == _T_90055 ? shiftedStoreDataQPreg_13 : _GEN_1766; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1768 = 4'he == _T_90055 ? shiftedStoreDataQPreg_14 : _GEN_1767; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign _GEN_1769 = 4'hf == _T_90055 ? shiftedStoreDataQPreg_15 : _GEN_1768; // @[AxiLoadQueue.scala 195:31:@36301.6]
  assign lastConflict_13_0 = _T_90072 ? _GEN_1722 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_1 = _T_90072 ? _GEN_1723 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_2 = _T_90072 ? _GEN_1724 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_3 = _T_90072 ? _GEN_1725 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_4 = _T_90072 ? _GEN_1726 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_5 = _T_90072 ? _GEN_1727 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_6 = _T_90072 ? _GEN_1728 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_7 = _T_90072 ? _GEN_1729 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_8 = _T_90072 ? _GEN_1730 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_9 = _T_90072 ? _GEN_1731 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_10 = _T_90072 ? _GEN_1732 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_11 = _T_90072 ? _GEN_1733 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_12 = _T_90072 ? _GEN_1734 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_13 = _T_90072 ? _GEN_1735 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_14 = _T_90072 ? _GEN_1736 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign lastConflict_13_15 = _T_90072 ? _GEN_1737 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign canBypass_13 = _T_90072 ? _GEN_1753 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign bypassVal_13 = _T_90072 ? _GEN_1769 : 32'h0; // @[AxiLoadQueue.scala 192:53:@36298.4]
  assign _T_90178 = conflictPReg_14_2 ? 2'h2 : {{1'd0}, conflictPReg_14_1}; // @[AxiLoadQueue.scala 191:60:@36355.4]
  assign _T_90179 = conflictPReg_14_3 ? 2'h3 : _T_90178; // @[AxiLoadQueue.scala 191:60:@36356.4]
  assign _T_90180 = conflictPReg_14_4 ? 3'h4 : {{1'd0}, _T_90179}; // @[AxiLoadQueue.scala 191:60:@36357.4]
  assign _T_90181 = conflictPReg_14_5 ? 3'h5 : _T_90180; // @[AxiLoadQueue.scala 191:60:@36358.4]
  assign _T_90182 = conflictPReg_14_6 ? 3'h6 : _T_90181; // @[AxiLoadQueue.scala 191:60:@36359.4]
  assign _T_90183 = conflictPReg_14_7 ? 3'h7 : _T_90182; // @[AxiLoadQueue.scala 191:60:@36360.4]
  assign _T_90184 = conflictPReg_14_8 ? 4'h8 : {{1'd0}, _T_90183}; // @[AxiLoadQueue.scala 191:60:@36361.4]
  assign _T_90185 = conflictPReg_14_9 ? 4'h9 : _T_90184; // @[AxiLoadQueue.scala 191:60:@36362.4]
  assign _T_90186 = conflictPReg_14_10 ? 4'ha : _T_90185; // @[AxiLoadQueue.scala 191:60:@36363.4]
  assign _T_90187 = conflictPReg_14_11 ? 4'hb : _T_90186; // @[AxiLoadQueue.scala 191:60:@36364.4]
  assign _T_90188 = conflictPReg_14_12 ? 4'hc : _T_90187; // @[AxiLoadQueue.scala 191:60:@36365.4]
  assign _T_90189 = conflictPReg_14_13 ? 4'hd : _T_90188; // @[AxiLoadQueue.scala 191:60:@36366.4]
  assign _T_90190 = conflictPReg_14_14 ? 4'he : _T_90189; // @[AxiLoadQueue.scala 191:60:@36367.4]
  assign _T_90191 = conflictPReg_14_15 ? 4'hf : _T_90190; // @[AxiLoadQueue.scala 191:60:@36368.4]
  assign _T_90194 = conflictPReg_14_0 | conflictPReg_14_1; // @[AxiLoadQueue.scala 192:43:@36370.4]
  assign _T_90195 = _T_90194 | conflictPReg_14_2; // @[AxiLoadQueue.scala 192:43:@36371.4]
  assign _T_90196 = _T_90195 | conflictPReg_14_3; // @[AxiLoadQueue.scala 192:43:@36372.4]
  assign _T_90197 = _T_90196 | conflictPReg_14_4; // @[AxiLoadQueue.scala 192:43:@36373.4]
  assign _T_90198 = _T_90197 | conflictPReg_14_5; // @[AxiLoadQueue.scala 192:43:@36374.4]
  assign _T_90199 = _T_90198 | conflictPReg_14_6; // @[AxiLoadQueue.scala 192:43:@36375.4]
  assign _T_90200 = _T_90199 | conflictPReg_14_7; // @[AxiLoadQueue.scala 192:43:@36376.4]
  assign _T_90201 = _T_90200 | conflictPReg_14_8; // @[AxiLoadQueue.scala 192:43:@36377.4]
  assign _T_90202 = _T_90201 | conflictPReg_14_9; // @[AxiLoadQueue.scala 192:43:@36378.4]
  assign _T_90203 = _T_90202 | conflictPReg_14_10; // @[AxiLoadQueue.scala 192:43:@36379.4]
  assign _T_90204 = _T_90203 | conflictPReg_14_11; // @[AxiLoadQueue.scala 192:43:@36380.4]
  assign _T_90205 = _T_90204 | conflictPReg_14_12; // @[AxiLoadQueue.scala 192:43:@36381.4]
  assign _T_90206 = _T_90205 | conflictPReg_14_13; // @[AxiLoadQueue.scala 192:43:@36382.4]
  assign _T_90207 = _T_90206 | conflictPReg_14_14; // @[AxiLoadQueue.scala 192:43:@36383.4]
  assign _T_90208 = _T_90207 | conflictPReg_14_15; // @[AxiLoadQueue.scala 192:43:@36384.4]
  assign _GEN_1788 = 4'h0 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1789 = 4'h1 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1790 = 4'h2 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1791 = 4'h3 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1792 = 4'h4 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1793 = 4'h5 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1794 = 4'h6 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1795 = 4'h7 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1796 = 4'h8 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1797 = 4'h9 == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1798 = 4'ha == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1799 = 4'hb == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1800 = 4'hc == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1801 = 4'hd == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1802 = 4'he == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1803 = 4'hf == _T_90191; // @[AxiLoadQueue.scala 193:43:@36386.6]
  assign _GEN_1805 = 4'h1 == _T_90191 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1806 = 4'h2 == _T_90191 ? shiftedStoreDataKnownPReg_2 : _GEN_1805; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1807 = 4'h3 == _T_90191 ? shiftedStoreDataKnownPReg_3 : _GEN_1806; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1808 = 4'h4 == _T_90191 ? shiftedStoreDataKnownPReg_4 : _GEN_1807; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1809 = 4'h5 == _T_90191 ? shiftedStoreDataKnownPReg_5 : _GEN_1808; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1810 = 4'h6 == _T_90191 ? shiftedStoreDataKnownPReg_6 : _GEN_1809; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1811 = 4'h7 == _T_90191 ? shiftedStoreDataKnownPReg_7 : _GEN_1810; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1812 = 4'h8 == _T_90191 ? shiftedStoreDataKnownPReg_8 : _GEN_1811; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1813 = 4'h9 == _T_90191 ? shiftedStoreDataKnownPReg_9 : _GEN_1812; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1814 = 4'ha == _T_90191 ? shiftedStoreDataKnownPReg_10 : _GEN_1813; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1815 = 4'hb == _T_90191 ? shiftedStoreDataKnownPReg_11 : _GEN_1814; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1816 = 4'hc == _T_90191 ? shiftedStoreDataKnownPReg_12 : _GEN_1815; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1817 = 4'hd == _T_90191 ? shiftedStoreDataKnownPReg_13 : _GEN_1816; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1818 = 4'he == _T_90191 ? shiftedStoreDataKnownPReg_14 : _GEN_1817; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1819 = 4'hf == _T_90191 ? shiftedStoreDataKnownPReg_15 : _GEN_1818; // @[AxiLoadQueue.scala 194:31:@36387.6]
  assign _GEN_1821 = 4'h1 == _T_90191 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1822 = 4'h2 == _T_90191 ? shiftedStoreDataQPreg_2 : _GEN_1821; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1823 = 4'h3 == _T_90191 ? shiftedStoreDataQPreg_3 : _GEN_1822; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1824 = 4'h4 == _T_90191 ? shiftedStoreDataQPreg_4 : _GEN_1823; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1825 = 4'h5 == _T_90191 ? shiftedStoreDataQPreg_5 : _GEN_1824; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1826 = 4'h6 == _T_90191 ? shiftedStoreDataQPreg_6 : _GEN_1825; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1827 = 4'h7 == _T_90191 ? shiftedStoreDataQPreg_7 : _GEN_1826; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1828 = 4'h8 == _T_90191 ? shiftedStoreDataQPreg_8 : _GEN_1827; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1829 = 4'h9 == _T_90191 ? shiftedStoreDataQPreg_9 : _GEN_1828; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1830 = 4'ha == _T_90191 ? shiftedStoreDataQPreg_10 : _GEN_1829; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1831 = 4'hb == _T_90191 ? shiftedStoreDataQPreg_11 : _GEN_1830; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1832 = 4'hc == _T_90191 ? shiftedStoreDataQPreg_12 : _GEN_1831; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1833 = 4'hd == _T_90191 ? shiftedStoreDataQPreg_13 : _GEN_1832; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1834 = 4'he == _T_90191 ? shiftedStoreDataQPreg_14 : _GEN_1833; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign _GEN_1835 = 4'hf == _T_90191 ? shiftedStoreDataQPreg_15 : _GEN_1834; // @[AxiLoadQueue.scala 195:31:@36388.6]
  assign lastConflict_14_0 = _T_90208 ? _GEN_1788 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_1 = _T_90208 ? _GEN_1789 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_2 = _T_90208 ? _GEN_1790 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_3 = _T_90208 ? _GEN_1791 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_4 = _T_90208 ? _GEN_1792 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_5 = _T_90208 ? _GEN_1793 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_6 = _T_90208 ? _GEN_1794 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_7 = _T_90208 ? _GEN_1795 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_8 = _T_90208 ? _GEN_1796 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_9 = _T_90208 ? _GEN_1797 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_10 = _T_90208 ? _GEN_1798 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_11 = _T_90208 ? _GEN_1799 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_12 = _T_90208 ? _GEN_1800 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_13 = _T_90208 ? _GEN_1801 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_14 = _T_90208 ? _GEN_1802 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign lastConflict_14_15 = _T_90208 ? _GEN_1803 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign canBypass_14 = _T_90208 ? _GEN_1819 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign bypassVal_14 = _T_90208 ? _GEN_1835 : 32'h0; // @[AxiLoadQueue.scala 192:53:@36385.4]
  assign _T_90314 = conflictPReg_15_2 ? 2'h2 : {{1'd0}, conflictPReg_15_1}; // @[AxiLoadQueue.scala 191:60:@36442.4]
  assign _T_90315 = conflictPReg_15_3 ? 2'h3 : _T_90314; // @[AxiLoadQueue.scala 191:60:@36443.4]
  assign _T_90316 = conflictPReg_15_4 ? 3'h4 : {{1'd0}, _T_90315}; // @[AxiLoadQueue.scala 191:60:@36444.4]
  assign _T_90317 = conflictPReg_15_5 ? 3'h5 : _T_90316; // @[AxiLoadQueue.scala 191:60:@36445.4]
  assign _T_90318 = conflictPReg_15_6 ? 3'h6 : _T_90317; // @[AxiLoadQueue.scala 191:60:@36446.4]
  assign _T_90319 = conflictPReg_15_7 ? 3'h7 : _T_90318; // @[AxiLoadQueue.scala 191:60:@36447.4]
  assign _T_90320 = conflictPReg_15_8 ? 4'h8 : {{1'd0}, _T_90319}; // @[AxiLoadQueue.scala 191:60:@36448.4]
  assign _T_90321 = conflictPReg_15_9 ? 4'h9 : _T_90320; // @[AxiLoadQueue.scala 191:60:@36449.4]
  assign _T_90322 = conflictPReg_15_10 ? 4'ha : _T_90321; // @[AxiLoadQueue.scala 191:60:@36450.4]
  assign _T_90323 = conflictPReg_15_11 ? 4'hb : _T_90322; // @[AxiLoadQueue.scala 191:60:@36451.4]
  assign _T_90324 = conflictPReg_15_12 ? 4'hc : _T_90323; // @[AxiLoadQueue.scala 191:60:@36452.4]
  assign _T_90325 = conflictPReg_15_13 ? 4'hd : _T_90324; // @[AxiLoadQueue.scala 191:60:@36453.4]
  assign _T_90326 = conflictPReg_15_14 ? 4'he : _T_90325; // @[AxiLoadQueue.scala 191:60:@36454.4]
  assign _T_90327 = conflictPReg_15_15 ? 4'hf : _T_90326; // @[AxiLoadQueue.scala 191:60:@36455.4]
  assign _T_90330 = conflictPReg_15_0 | conflictPReg_15_1; // @[AxiLoadQueue.scala 192:43:@36457.4]
  assign _T_90331 = _T_90330 | conflictPReg_15_2; // @[AxiLoadQueue.scala 192:43:@36458.4]
  assign _T_90332 = _T_90331 | conflictPReg_15_3; // @[AxiLoadQueue.scala 192:43:@36459.4]
  assign _T_90333 = _T_90332 | conflictPReg_15_4; // @[AxiLoadQueue.scala 192:43:@36460.4]
  assign _T_90334 = _T_90333 | conflictPReg_15_5; // @[AxiLoadQueue.scala 192:43:@36461.4]
  assign _T_90335 = _T_90334 | conflictPReg_15_6; // @[AxiLoadQueue.scala 192:43:@36462.4]
  assign _T_90336 = _T_90335 | conflictPReg_15_7; // @[AxiLoadQueue.scala 192:43:@36463.4]
  assign _T_90337 = _T_90336 | conflictPReg_15_8; // @[AxiLoadQueue.scala 192:43:@36464.4]
  assign _T_90338 = _T_90337 | conflictPReg_15_9; // @[AxiLoadQueue.scala 192:43:@36465.4]
  assign _T_90339 = _T_90338 | conflictPReg_15_10; // @[AxiLoadQueue.scala 192:43:@36466.4]
  assign _T_90340 = _T_90339 | conflictPReg_15_11; // @[AxiLoadQueue.scala 192:43:@36467.4]
  assign _T_90341 = _T_90340 | conflictPReg_15_12; // @[AxiLoadQueue.scala 192:43:@36468.4]
  assign _T_90342 = _T_90341 | conflictPReg_15_13; // @[AxiLoadQueue.scala 192:43:@36469.4]
  assign _T_90343 = _T_90342 | conflictPReg_15_14; // @[AxiLoadQueue.scala 192:43:@36470.4]
  assign _T_90344 = _T_90343 | conflictPReg_15_15; // @[AxiLoadQueue.scala 192:43:@36471.4]
  assign _GEN_1854 = 4'h0 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1855 = 4'h1 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1856 = 4'h2 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1857 = 4'h3 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1858 = 4'h4 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1859 = 4'h5 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1860 = 4'h6 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1861 = 4'h7 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1862 = 4'h8 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1863 = 4'h9 == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1864 = 4'ha == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1865 = 4'hb == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1866 = 4'hc == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1867 = 4'hd == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1868 = 4'he == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1869 = 4'hf == _T_90327; // @[AxiLoadQueue.scala 193:43:@36473.6]
  assign _GEN_1871 = 4'h1 == _T_90327 ? shiftedStoreDataKnownPReg_1 : shiftedStoreDataKnownPReg_0; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1872 = 4'h2 == _T_90327 ? shiftedStoreDataKnownPReg_2 : _GEN_1871; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1873 = 4'h3 == _T_90327 ? shiftedStoreDataKnownPReg_3 : _GEN_1872; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1874 = 4'h4 == _T_90327 ? shiftedStoreDataKnownPReg_4 : _GEN_1873; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1875 = 4'h5 == _T_90327 ? shiftedStoreDataKnownPReg_5 : _GEN_1874; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1876 = 4'h6 == _T_90327 ? shiftedStoreDataKnownPReg_6 : _GEN_1875; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1877 = 4'h7 == _T_90327 ? shiftedStoreDataKnownPReg_7 : _GEN_1876; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1878 = 4'h8 == _T_90327 ? shiftedStoreDataKnownPReg_8 : _GEN_1877; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1879 = 4'h9 == _T_90327 ? shiftedStoreDataKnownPReg_9 : _GEN_1878; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1880 = 4'ha == _T_90327 ? shiftedStoreDataKnownPReg_10 : _GEN_1879; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1881 = 4'hb == _T_90327 ? shiftedStoreDataKnownPReg_11 : _GEN_1880; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1882 = 4'hc == _T_90327 ? shiftedStoreDataKnownPReg_12 : _GEN_1881; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1883 = 4'hd == _T_90327 ? shiftedStoreDataKnownPReg_13 : _GEN_1882; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1884 = 4'he == _T_90327 ? shiftedStoreDataKnownPReg_14 : _GEN_1883; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1885 = 4'hf == _T_90327 ? shiftedStoreDataKnownPReg_15 : _GEN_1884; // @[AxiLoadQueue.scala 194:31:@36474.6]
  assign _GEN_1887 = 4'h1 == _T_90327 ? shiftedStoreDataQPreg_1 : shiftedStoreDataQPreg_0; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1888 = 4'h2 == _T_90327 ? shiftedStoreDataQPreg_2 : _GEN_1887; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1889 = 4'h3 == _T_90327 ? shiftedStoreDataQPreg_3 : _GEN_1888; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1890 = 4'h4 == _T_90327 ? shiftedStoreDataQPreg_4 : _GEN_1889; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1891 = 4'h5 == _T_90327 ? shiftedStoreDataQPreg_5 : _GEN_1890; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1892 = 4'h6 == _T_90327 ? shiftedStoreDataQPreg_6 : _GEN_1891; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1893 = 4'h7 == _T_90327 ? shiftedStoreDataQPreg_7 : _GEN_1892; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1894 = 4'h8 == _T_90327 ? shiftedStoreDataQPreg_8 : _GEN_1893; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1895 = 4'h9 == _T_90327 ? shiftedStoreDataQPreg_9 : _GEN_1894; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1896 = 4'ha == _T_90327 ? shiftedStoreDataQPreg_10 : _GEN_1895; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1897 = 4'hb == _T_90327 ? shiftedStoreDataQPreg_11 : _GEN_1896; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1898 = 4'hc == _T_90327 ? shiftedStoreDataQPreg_12 : _GEN_1897; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1899 = 4'hd == _T_90327 ? shiftedStoreDataQPreg_13 : _GEN_1898; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1900 = 4'he == _T_90327 ? shiftedStoreDataQPreg_14 : _GEN_1899; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign _GEN_1901 = 4'hf == _T_90327 ? shiftedStoreDataQPreg_15 : _GEN_1900; // @[AxiLoadQueue.scala 195:31:@36475.6]
  assign lastConflict_15_0 = _T_90344 ? _GEN_1854 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_1 = _T_90344 ? _GEN_1855 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_2 = _T_90344 ? _GEN_1856 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_3 = _T_90344 ? _GEN_1857 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_4 = _T_90344 ? _GEN_1858 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_5 = _T_90344 ? _GEN_1859 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_6 = _T_90344 ? _GEN_1860 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_7 = _T_90344 ? _GEN_1861 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_8 = _T_90344 ? _GEN_1862 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_9 = _T_90344 ? _GEN_1863 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_10 = _T_90344 ? _GEN_1864 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_11 = _T_90344 ? _GEN_1865 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_12 = _T_90344 ? _GEN_1866 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_13 = _T_90344 ? _GEN_1867 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_14 = _T_90344 ? _GEN_1868 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign lastConflict_15_15 = _T_90344 ? _GEN_1869 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign canBypass_15 = _T_90344 ? _GEN_1885 : 1'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign bypassVal_15 = _T_90344 ? _GEN_1901 : 32'h0; // @[AxiLoadQueue.scala 192:53:@36472.4]
  assign _T_90404 = 16'h1 << head; // @[OneHot.scala 52:12:@36480.4]
  assign _T_90406 = _T_90404[0]; // @[util.scala 33:60:@36482.4]
  assign _T_90407 = _T_90404[1]; // @[util.scala 33:60:@36483.4]
  assign _T_90408 = _T_90404[2]; // @[util.scala 33:60:@36484.4]
  assign _T_90409 = _T_90404[3]; // @[util.scala 33:60:@36485.4]
  assign _T_90410 = _T_90404[4]; // @[util.scala 33:60:@36486.4]
  assign _T_90411 = _T_90404[5]; // @[util.scala 33:60:@36487.4]
  assign _T_90412 = _T_90404[6]; // @[util.scala 33:60:@36488.4]
  assign _T_90413 = _T_90404[7]; // @[util.scala 33:60:@36489.4]
  assign _T_90414 = _T_90404[8]; // @[util.scala 33:60:@36490.4]
  assign _T_90415 = _T_90404[9]; // @[util.scala 33:60:@36491.4]
  assign _T_90416 = _T_90404[10]; // @[util.scala 33:60:@36492.4]
  assign _T_90417 = _T_90404[11]; // @[util.scala 33:60:@36493.4]
  assign _T_90418 = _T_90404[12]; // @[util.scala 33:60:@36494.4]
  assign _T_90419 = _T_90404[13]; // @[util.scala 33:60:@36495.4]
  assign _T_90420 = _T_90404[14]; // @[util.scala 33:60:@36496.4]
  assign _T_90421 = _T_90404[15]; // @[util.scala 33:60:@36497.4]
  assign _T_93610 = dataKnownPReg_15 == 1'h0; // @[AxiLoadQueue.scala 242:41:@39144.4]
  assign _T_93611 = addrKnownPReg_15 & _T_93610; // @[AxiLoadQueue.scala 242:38:@39145.4]
  assign _T_93613 = bypassInitiated_15 == 1'h0; // @[AxiLoadQueue.scala 243:12:@39147.6]
  assign _T_93615 = loadInitiated_15 == 1'h0; // @[AxiLoadQueue.scala 243:46:@39148.6]
  assign _T_93616 = _T_93613 & _T_93615; // @[AxiLoadQueue.scala 243:43:@39149.6]
  assign _T_93618 = dataKnown_15 == 1'h0; // @[AxiLoadQueue.scala 243:78:@39150.6]
  assign _T_93619 = _T_93616 & _T_93618; // @[AxiLoadQueue.scala 243:75:@39151.6]
  assign _T_93622 = storeAddrNotKnownFlagsPReg_15_0 | storeAddrNotKnownFlagsPReg_15_1; // @[AxiLoadQueue.scala 246:86:@39154.8]
  assign _T_93623 = _T_93622 | storeAddrNotKnownFlagsPReg_15_2; // @[AxiLoadQueue.scala 246:86:@39155.8]
  assign _T_93624 = _T_93623 | storeAddrNotKnownFlagsPReg_15_3; // @[AxiLoadQueue.scala 246:86:@39156.8]
  assign _T_93625 = _T_93624 | storeAddrNotKnownFlagsPReg_15_4; // @[AxiLoadQueue.scala 246:86:@39157.8]
  assign _T_93626 = _T_93625 | storeAddrNotKnownFlagsPReg_15_5; // @[AxiLoadQueue.scala 246:86:@39158.8]
  assign _T_93627 = _T_93626 | storeAddrNotKnownFlagsPReg_15_6; // @[AxiLoadQueue.scala 246:86:@39159.8]
  assign _T_93628 = _T_93627 | storeAddrNotKnownFlagsPReg_15_7; // @[AxiLoadQueue.scala 246:86:@39160.8]
  assign _T_93629 = _T_93628 | storeAddrNotKnownFlagsPReg_15_8; // @[AxiLoadQueue.scala 246:86:@39161.8]
  assign _T_93630 = _T_93629 | storeAddrNotKnownFlagsPReg_15_9; // @[AxiLoadQueue.scala 246:86:@39162.8]
  assign _T_93631 = _T_93630 | storeAddrNotKnownFlagsPReg_15_10; // @[AxiLoadQueue.scala 246:86:@39163.8]
  assign _T_93632 = _T_93631 | storeAddrNotKnownFlagsPReg_15_11; // @[AxiLoadQueue.scala 246:86:@39164.8]
  assign _T_93633 = _T_93632 | storeAddrNotKnownFlagsPReg_15_12; // @[AxiLoadQueue.scala 246:86:@39165.8]
  assign _T_93634 = _T_93633 | storeAddrNotKnownFlagsPReg_15_13; // @[AxiLoadQueue.scala 246:86:@39166.8]
  assign _T_93635 = _T_93634 | storeAddrNotKnownFlagsPReg_15_14; // @[AxiLoadQueue.scala 246:86:@39167.8]
  assign _T_93636 = _T_93635 | storeAddrNotKnownFlagsPReg_15_15; // @[AxiLoadQueue.scala 246:86:@39168.8]
  assign _T_93638 = _T_93636 == 1'h0; // @[AxiLoadQueue.scala 246:38:@39169.8]
  assign _T_93657 = _T_90344 == 1'h0; // @[AxiLoadQueue.scala 247:11:@39186.8]
  assign _T_93658 = _T_93638 & _T_93657; // @[AxiLoadQueue.scala 246:103:@39187.8]
  assign _GEN_2060 = _T_93619 ? _T_93658 : 1'h0; // @[AxiLoadQueue.scala 243:104:@39152.6]
  assign loadRequest_15 = _T_93611 ? _GEN_2060 : 1'h0; // @[AxiLoadQueue.scala 242:71:@39146.4]
  assign _T_90462 = loadRequest_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36515.4]
  assign _T_93526 = dataKnownPReg_14 == 1'h0; // @[AxiLoadQueue.scala 242:41:@39062.4]
  assign _T_93527 = addrKnownPReg_14 & _T_93526; // @[AxiLoadQueue.scala 242:38:@39063.4]
  assign _T_93529 = bypassInitiated_14 == 1'h0; // @[AxiLoadQueue.scala 243:12:@39065.6]
  assign _T_93531 = loadInitiated_14 == 1'h0; // @[AxiLoadQueue.scala 243:46:@39066.6]
  assign _T_93532 = _T_93529 & _T_93531; // @[AxiLoadQueue.scala 243:43:@39067.6]
  assign _T_93534 = dataKnown_14 == 1'h0; // @[AxiLoadQueue.scala 243:78:@39068.6]
  assign _T_93535 = _T_93532 & _T_93534; // @[AxiLoadQueue.scala 243:75:@39069.6]
  assign _T_93538 = storeAddrNotKnownFlagsPReg_14_0 | storeAddrNotKnownFlagsPReg_14_1; // @[AxiLoadQueue.scala 246:86:@39072.8]
  assign _T_93539 = _T_93538 | storeAddrNotKnownFlagsPReg_14_2; // @[AxiLoadQueue.scala 246:86:@39073.8]
  assign _T_93540 = _T_93539 | storeAddrNotKnownFlagsPReg_14_3; // @[AxiLoadQueue.scala 246:86:@39074.8]
  assign _T_93541 = _T_93540 | storeAddrNotKnownFlagsPReg_14_4; // @[AxiLoadQueue.scala 246:86:@39075.8]
  assign _T_93542 = _T_93541 | storeAddrNotKnownFlagsPReg_14_5; // @[AxiLoadQueue.scala 246:86:@39076.8]
  assign _T_93543 = _T_93542 | storeAddrNotKnownFlagsPReg_14_6; // @[AxiLoadQueue.scala 246:86:@39077.8]
  assign _T_93544 = _T_93543 | storeAddrNotKnownFlagsPReg_14_7; // @[AxiLoadQueue.scala 246:86:@39078.8]
  assign _T_93545 = _T_93544 | storeAddrNotKnownFlagsPReg_14_8; // @[AxiLoadQueue.scala 246:86:@39079.8]
  assign _T_93546 = _T_93545 | storeAddrNotKnownFlagsPReg_14_9; // @[AxiLoadQueue.scala 246:86:@39080.8]
  assign _T_93547 = _T_93546 | storeAddrNotKnownFlagsPReg_14_10; // @[AxiLoadQueue.scala 246:86:@39081.8]
  assign _T_93548 = _T_93547 | storeAddrNotKnownFlagsPReg_14_11; // @[AxiLoadQueue.scala 246:86:@39082.8]
  assign _T_93549 = _T_93548 | storeAddrNotKnownFlagsPReg_14_12; // @[AxiLoadQueue.scala 246:86:@39083.8]
  assign _T_93550 = _T_93549 | storeAddrNotKnownFlagsPReg_14_13; // @[AxiLoadQueue.scala 246:86:@39084.8]
  assign _T_93551 = _T_93550 | storeAddrNotKnownFlagsPReg_14_14; // @[AxiLoadQueue.scala 246:86:@39085.8]
  assign _T_93552 = _T_93551 | storeAddrNotKnownFlagsPReg_14_15; // @[AxiLoadQueue.scala 246:86:@39086.8]
  assign _T_93554 = _T_93552 == 1'h0; // @[AxiLoadQueue.scala 246:38:@39087.8]
  assign _T_93573 = _T_90208 == 1'h0; // @[AxiLoadQueue.scala 247:11:@39104.8]
  assign _T_93574 = _T_93554 & _T_93573; // @[AxiLoadQueue.scala 246:103:@39105.8]
  assign _GEN_2056 = _T_93535 ? _T_93574 : 1'h0; // @[AxiLoadQueue.scala 243:104:@39070.6]
  assign loadRequest_14 = _T_93527 ? _GEN_2056 : 1'h0; // @[AxiLoadQueue.scala 242:71:@39064.4]
  assign _T_90463 = loadRequest_14 ? 16'h4000 : _T_90462; // @[Mux.scala 31:69:@36516.4]
  assign _T_93442 = dataKnownPReg_13 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38980.4]
  assign _T_93443 = addrKnownPReg_13 & _T_93442; // @[AxiLoadQueue.scala 242:38:@38981.4]
  assign _T_93445 = bypassInitiated_13 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38983.6]
  assign _T_93447 = loadInitiated_13 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38984.6]
  assign _T_93448 = _T_93445 & _T_93447; // @[AxiLoadQueue.scala 243:43:@38985.6]
  assign _T_93450 = dataKnown_13 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38986.6]
  assign _T_93451 = _T_93448 & _T_93450; // @[AxiLoadQueue.scala 243:75:@38987.6]
  assign _T_93454 = storeAddrNotKnownFlagsPReg_13_0 | storeAddrNotKnownFlagsPReg_13_1; // @[AxiLoadQueue.scala 246:86:@38990.8]
  assign _T_93455 = _T_93454 | storeAddrNotKnownFlagsPReg_13_2; // @[AxiLoadQueue.scala 246:86:@38991.8]
  assign _T_93456 = _T_93455 | storeAddrNotKnownFlagsPReg_13_3; // @[AxiLoadQueue.scala 246:86:@38992.8]
  assign _T_93457 = _T_93456 | storeAddrNotKnownFlagsPReg_13_4; // @[AxiLoadQueue.scala 246:86:@38993.8]
  assign _T_93458 = _T_93457 | storeAddrNotKnownFlagsPReg_13_5; // @[AxiLoadQueue.scala 246:86:@38994.8]
  assign _T_93459 = _T_93458 | storeAddrNotKnownFlagsPReg_13_6; // @[AxiLoadQueue.scala 246:86:@38995.8]
  assign _T_93460 = _T_93459 | storeAddrNotKnownFlagsPReg_13_7; // @[AxiLoadQueue.scala 246:86:@38996.8]
  assign _T_93461 = _T_93460 | storeAddrNotKnownFlagsPReg_13_8; // @[AxiLoadQueue.scala 246:86:@38997.8]
  assign _T_93462 = _T_93461 | storeAddrNotKnownFlagsPReg_13_9; // @[AxiLoadQueue.scala 246:86:@38998.8]
  assign _T_93463 = _T_93462 | storeAddrNotKnownFlagsPReg_13_10; // @[AxiLoadQueue.scala 246:86:@38999.8]
  assign _T_93464 = _T_93463 | storeAddrNotKnownFlagsPReg_13_11; // @[AxiLoadQueue.scala 246:86:@39000.8]
  assign _T_93465 = _T_93464 | storeAddrNotKnownFlagsPReg_13_12; // @[AxiLoadQueue.scala 246:86:@39001.8]
  assign _T_93466 = _T_93465 | storeAddrNotKnownFlagsPReg_13_13; // @[AxiLoadQueue.scala 246:86:@39002.8]
  assign _T_93467 = _T_93466 | storeAddrNotKnownFlagsPReg_13_14; // @[AxiLoadQueue.scala 246:86:@39003.8]
  assign _T_93468 = _T_93467 | storeAddrNotKnownFlagsPReg_13_15; // @[AxiLoadQueue.scala 246:86:@39004.8]
  assign _T_93470 = _T_93468 == 1'h0; // @[AxiLoadQueue.scala 246:38:@39005.8]
  assign _T_93489 = _T_90072 == 1'h0; // @[AxiLoadQueue.scala 247:11:@39022.8]
  assign _T_93490 = _T_93470 & _T_93489; // @[AxiLoadQueue.scala 246:103:@39023.8]
  assign _GEN_2052 = _T_93451 ? _T_93490 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38988.6]
  assign loadRequest_13 = _T_93443 ? _GEN_2052 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38982.4]
  assign _T_90464 = loadRequest_13 ? 16'h2000 : _T_90463; // @[Mux.scala 31:69:@36517.4]
  assign _T_93358 = dataKnownPReg_12 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38898.4]
  assign _T_93359 = addrKnownPReg_12 & _T_93358; // @[AxiLoadQueue.scala 242:38:@38899.4]
  assign _T_93361 = bypassInitiated_12 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38901.6]
  assign _T_93363 = loadInitiated_12 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38902.6]
  assign _T_93364 = _T_93361 & _T_93363; // @[AxiLoadQueue.scala 243:43:@38903.6]
  assign _T_93366 = dataKnown_12 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38904.6]
  assign _T_93367 = _T_93364 & _T_93366; // @[AxiLoadQueue.scala 243:75:@38905.6]
  assign _T_93370 = storeAddrNotKnownFlagsPReg_12_0 | storeAddrNotKnownFlagsPReg_12_1; // @[AxiLoadQueue.scala 246:86:@38908.8]
  assign _T_93371 = _T_93370 | storeAddrNotKnownFlagsPReg_12_2; // @[AxiLoadQueue.scala 246:86:@38909.8]
  assign _T_93372 = _T_93371 | storeAddrNotKnownFlagsPReg_12_3; // @[AxiLoadQueue.scala 246:86:@38910.8]
  assign _T_93373 = _T_93372 | storeAddrNotKnownFlagsPReg_12_4; // @[AxiLoadQueue.scala 246:86:@38911.8]
  assign _T_93374 = _T_93373 | storeAddrNotKnownFlagsPReg_12_5; // @[AxiLoadQueue.scala 246:86:@38912.8]
  assign _T_93375 = _T_93374 | storeAddrNotKnownFlagsPReg_12_6; // @[AxiLoadQueue.scala 246:86:@38913.8]
  assign _T_93376 = _T_93375 | storeAddrNotKnownFlagsPReg_12_7; // @[AxiLoadQueue.scala 246:86:@38914.8]
  assign _T_93377 = _T_93376 | storeAddrNotKnownFlagsPReg_12_8; // @[AxiLoadQueue.scala 246:86:@38915.8]
  assign _T_93378 = _T_93377 | storeAddrNotKnownFlagsPReg_12_9; // @[AxiLoadQueue.scala 246:86:@38916.8]
  assign _T_93379 = _T_93378 | storeAddrNotKnownFlagsPReg_12_10; // @[AxiLoadQueue.scala 246:86:@38917.8]
  assign _T_93380 = _T_93379 | storeAddrNotKnownFlagsPReg_12_11; // @[AxiLoadQueue.scala 246:86:@38918.8]
  assign _T_93381 = _T_93380 | storeAddrNotKnownFlagsPReg_12_12; // @[AxiLoadQueue.scala 246:86:@38919.8]
  assign _T_93382 = _T_93381 | storeAddrNotKnownFlagsPReg_12_13; // @[AxiLoadQueue.scala 246:86:@38920.8]
  assign _T_93383 = _T_93382 | storeAddrNotKnownFlagsPReg_12_14; // @[AxiLoadQueue.scala 246:86:@38921.8]
  assign _T_93384 = _T_93383 | storeAddrNotKnownFlagsPReg_12_15; // @[AxiLoadQueue.scala 246:86:@38922.8]
  assign _T_93386 = _T_93384 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38923.8]
  assign _T_93405 = _T_89936 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38940.8]
  assign _T_93406 = _T_93386 & _T_93405; // @[AxiLoadQueue.scala 246:103:@38941.8]
  assign _GEN_2048 = _T_93367 ? _T_93406 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38906.6]
  assign loadRequest_12 = _T_93359 ? _GEN_2048 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38900.4]
  assign _T_90465 = loadRequest_12 ? 16'h1000 : _T_90464; // @[Mux.scala 31:69:@36518.4]
  assign _T_93274 = dataKnownPReg_11 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38816.4]
  assign _T_93275 = addrKnownPReg_11 & _T_93274; // @[AxiLoadQueue.scala 242:38:@38817.4]
  assign _T_93277 = bypassInitiated_11 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38819.6]
  assign _T_93279 = loadInitiated_11 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38820.6]
  assign _T_93280 = _T_93277 & _T_93279; // @[AxiLoadQueue.scala 243:43:@38821.6]
  assign _T_93282 = dataKnown_11 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38822.6]
  assign _T_93283 = _T_93280 & _T_93282; // @[AxiLoadQueue.scala 243:75:@38823.6]
  assign _T_93286 = storeAddrNotKnownFlagsPReg_11_0 | storeAddrNotKnownFlagsPReg_11_1; // @[AxiLoadQueue.scala 246:86:@38826.8]
  assign _T_93287 = _T_93286 | storeAddrNotKnownFlagsPReg_11_2; // @[AxiLoadQueue.scala 246:86:@38827.8]
  assign _T_93288 = _T_93287 | storeAddrNotKnownFlagsPReg_11_3; // @[AxiLoadQueue.scala 246:86:@38828.8]
  assign _T_93289 = _T_93288 | storeAddrNotKnownFlagsPReg_11_4; // @[AxiLoadQueue.scala 246:86:@38829.8]
  assign _T_93290 = _T_93289 | storeAddrNotKnownFlagsPReg_11_5; // @[AxiLoadQueue.scala 246:86:@38830.8]
  assign _T_93291 = _T_93290 | storeAddrNotKnownFlagsPReg_11_6; // @[AxiLoadQueue.scala 246:86:@38831.8]
  assign _T_93292 = _T_93291 | storeAddrNotKnownFlagsPReg_11_7; // @[AxiLoadQueue.scala 246:86:@38832.8]
  assign _T_93293 = _T_93292 | storeAddrNotKnownFlagsPReg_11_8; // @[AxiLoadQueue.scala 246:86:@38833.8]
  assign _T_93294 = _T_93293 | storeAddrNotKnownFlagsPReg_11_9; // @[AxiLoadQueue.scala 246:86:@38834.8]
  assign _T_93295 = _T_93294 | storeAddrNotKnownFlagsPReg_11_10; // @[AxiLoadQueue.scala 246:86:@38835.8]
  assign _T_93296 = _T_93295 | storeAddrNotKnownFlagsPReg_11_11; // @[AxiLoadQueue.scala 246:86:@38836.8]
  assign _T_93297 = _T_93296 | storeAddrNotKnownFlagsPReg_11_12; // @[AxiLoadQueue.scala 246:86:@38837.8]
  assign _T_93298 = _T_93297 | storeAddrNotKnownFlagsPReg_11_13; // @[AxiLoadQueue.scala 246:86:@38838.8]
  assign _T_93299 = _T_93298 | storeAddrNotKnownFlagsPReg_11_14; // @[AxiLoadQueue.scala 246:86:@38839.8]
  assign _T_93300 = _T_93299 | storeAddrNotKnownFlagsPReg_11_15; // @[AxiLoadQueue.scala 246:86:@38840.8]
  assign _T_93302 = _T_93300 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38841.8]
  assign _T_93321 = _T_89800 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38858.8]
  assign _T_93322 = _T_93302 & _T_93321; // @[AxiLoadQueue.scala 246:103:@38859.8]
  assign _GEN_2044 = _T_93283 ? _T_93322 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38824.6]
  assign loadRequest_11 = _T_93275 ? _GEN_2044 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38818.4]
  assign _T_90466 = loadRequest_11 ? 16'h800 : _T_90465; // @[Mux.scala 31:69:@36519.4]
  assign _T_93190 = dataKnownPReg_10 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38734.4]
  assign _T_93191 = addrKnownPReg_10 & _T_93190; // @[AxiLoadQueue.scala 242:38:@38735.4]
  assign _T_93193 = bypassInitiated_10 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38737.6]
  assign _T_93195 = loadInitiated_10 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38738.6]
  assign _T_93196 = _T_93193 & _T_93195; // @[AxiLoadQueue.scala 243:43:@38739.6]
  assign _T_93198 = dataKnown_10 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38740.6]
  assign _T_93199 = _T_93196 & _T_93198; // @[AxiLoadQueue.scala 243:75:@38741.6]
  assign _T_93202 = storeAddrNotKnownFlagsPReg_10_0 | storeAddrNotKnownFlagsPReg_10_1; // @[AxiLoadQueue.scala 246:86:@38744.8]
  assign _T_93203 = _T_93202 | storeAddrNotKnownFlagsPReg_10_2; // @[AxiLoadQueue.scala 246:86:@38745.8]
  assign _T_93204 = _T_93203 | storeAddrNotKnownFlagsPReg_10_3; // @[AxiLoadQueue.scala 246:86:@38746.8]
  assign _T_93205 = _T_93204 | storeAddrNotKnownFlagsPReg_10_4; // @[AxiLoadQueue.scala 246:86:@38747.8]
  assign _T_93206 = _T_93205 | storeAddrNotKnownFlagsPReg_10_5; // @[AxiLoadQueue.scala 246:86:@38748.8]
  assign _T_93207 = _T_93206 | storeAddrNotKnownFlagsPReg_10_6; // @[AxiLoadQueue.scala 246:86:@38749.8]
  assign _T_93208 = _T_93207 | storeAddrNotKnownFlagsPReg_10_7; // @[AxiLoadQueue.scala 246:86:@38750.8]
  assign _T_93209 = _T_93208 | storeAddrNotKnownFlagsPReg_10_8; // @[AxiLoadQueue.scala 246:86:@38751.8]
  assign _T_93210 = _T_93209 | storeAddrNotKnownFlagsPReg_10_9; // @[AxiLoadQueue.scala 246:86:@38752.8]
  assign _T_93211 = _T_93210 | storeAddrNotKnownFlagsPReg_10_10; // @[AxiLoadQueue.scala 246:86:@38753.8]
  assign _T_93212 = _T_93211 | storeAddrNotKnownFlagsPReg_10_11; // @[AxiLoadQueue.scala 246:86:@38754.8]
  assign _T_93213 = _T_93212 | storeAddrNotKnownFlagsPReg_10_12; // @[AxiLoadQueue.scala 246:86:@38755.8]
  assign _T_93214 = _T_93213 | storeAddrNotKnownFlagsPReg_10_13; // @[AxiLoadQueue.scala 246:86:@38756.8]
  assign _T_93215 = _T_93214 | storeAddrNotKnownFlagsPReg_10_14; // @[AxiLoadQueue.scala 246:86:@38757.8]
  assign _T_93216 = _T_93215 | storeAddrNotKnownFlagsPReg_10_15; // @[AxiLoadQueue.scala 246:86:@38758.8]
  assign _T_93218 = _T_93216 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38759.8]
  assign _T_93237 = _T_89664 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38776.8]
  assign _T_93238 = _T_93218 & _T_93237; // @[AxiLoadQueue.scala 246:103:@38777.8]
  assign _GEN_2040 = _T_93199 ? _T_93238 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38742.6]
  assign loadRequest_10 = _T_93191 ? _GEN_2040 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38736.4]
  assign _T_90467 = loadRequest_10 ? 16'h400 : _T_90466; // @[Mux.scala 31:69:@36520.4]
  assign _T_93106 = dataKnownPReg_9 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38652.4]
  assign _T_93107 = addrKnownPReg_9 & _T_93106; // @[AxiLoadQueue.scala 242:38:@38653.4]
  assign _T_93109 = bypassInitiated_9 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38655.6]
  assign _T_93111 = loadInitiated_9 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38656.6]
  assign _T_93112 = _T_93109 & _T_93111; // @[AxiLoadQueue.scala 243:43:@38657.6]
  assign _T_93114 = dataKnown_9 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38658.6]
  assign _T_93115 = _T_93112 & _T_93114; // @[AxiLoadQueue.scala 243:75:@38659.6]
  assign _T_93118 = storeAddrNotKnownFlagsPReg_9_0 | storeAddrNotKnownFlagsPReg_9_1; // @[AxiLoadQueue.scala 246:86:@38662.8]
  assign _T_93119 = _T_93118 | storeAddrNotKnownFlagsPReg_9_2; // @[AxiLoadQueue.scala 246:86:@38663.8]
  assign _T_93120 = _T_93119 | storeAddrNotKnownFlagsPReg_9_3; // @[AxiLoadQueue.scala 246:86:@38664.8]
  assign _T_93121 = _T_93120 | storeAddrNotKnownFlagsPReg_9_4; // @[AxiLoadQueue.scala 246:86:@38665.8]
  assign _T_93122 = _T_93121 | storeAddrNotKnownFlagsPReg_9_5; // @[AxiLoadQueue.scala 246:86:@38666.8]
  assign _T_93123 = _T_93122 | storeAddrNotKnownFlagsPReg_9_6; // @[AxiLoadQueue.scala 246:86:@38667.8]
  assign _T_93124 = _T_93123 | storeAddrNotKnownFlagsPReg_9_7; // @[AxiLoadQueue.scala 246:86:@38668.8]
  assign _T_93125 = _T_93124 | storeAddrNotKnownFlagsPReg_9_8; // @[AxiLoadQueue.scala 246:86:@38669.8]
  assign _T_93126 = _T_93125 | storeAddrNotKnownFlagsPReg_9_9; // @[AxiLoadQueue.scala 246:86:@38670.8]
  assign _T_93127 = _T_93126 | storeAddrNotKnownFlagsPReg_9_10; // @[AxiLoadQueue.scala 246:86:@38671.8]
  assign _T_93128 = _T_93127 | storeAddrNotKnownFlagsPReg_9_11; // @[AxiLoadQueue.scala 246:86:@38672.8]
  assign _T_93129 = _T_93128 | storeAddrNotKnownFlagsPReg_9_12; // @[AxiLoadQueue.scala 246:86:@38673.8]
  assign _T_93130 = _T_93129 | storeAddrNotKnownFlagsPReg_9_13; // @[AxiLoadQueue.scala 246:86:@38674.8]
  assign _T_93131 = _T_93130 | storeAddrNotKnownFlagsPReg_9_14; // @[AxiLoadQueue.scala 246:86:@38675.8]
  assign _T_93132 = _T_93131 | storeAddrNotKnownFlagsPReg_9_15; // @[AxiLoadQueue.scala 246:86:@38676.8]
  assign _T_93134 = _T_93132 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38677.8]
  assign _T_93153 = _T_89528 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38694.8]
  assign _T_93154 = _T_93134 & _T_93153; // @[AxiLoadQueue.scala 246:103:@38695.8]
  assign _GEN_2036 = _T_93115 ? _T_93154 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38660.6]
  assign loadRequest_9 = _T_93107 ? _GEN_2036 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38654.4]
  assign _T_90468 = loadRequest_9 ? 16'h200 : _T_90467; // @[Mux.scala 31:69:@36521.4]
  assign _T_93022 = dataKnownPReg_8 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38570.4]
  assign _T_93023 = addrKnownPReg_8 & _T_93022; // @[AxiLoadQueue.scala 242:38:@38571.4]
  assign _T_93025 = bypassInitiated_8 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38573.6]
  assign _T_93027 = loadInitiated_8 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38574.6]
  assign _T_93028 = _T_93025 & _T_93027; // @[AxiLoadQueue.scala 243:43:@38575.6]
  assign _T_93030 = dataKnown_8 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38576.6]
  assign _T_93031 = _T_93028 & _T_93030; // @[AxiLoadQueue.scala 243:75:@38577.6]
  assign _T_93034 = storeAddrNotKnownFlagsPReg_8_0 | storeAddrNotKnownFlagsPReg_8_1; // @[AxiLoadQueue.scala 246:86:@38580.8]
  assign _T_93035 = _T_93034 | storeAddrNotKnownFlagsPReg_8_2; // @[AxiLoadQueue.scala 246:86:@38581.8]
  assign _T_93036 = _T_93035 | storeAddrNotKnownFlagsPReg_8_3; // @[AxiLoadQueue.scala 246:86:@38582.8]
  assign _T_93037 = _T_93036 | storeAddrNotKnownFlagsPReg_8_4; // @[AxiLoadQueue.scala 246:86:@38583.8]
  assign _T_93038 = _T_93037 | storeAddrNotKnownFlagsPReg_8_5; // @[AxiLoadQueue.scala 246:86:@38584.8]
  assign _T_93039 = _T_93038 | storeAddrNotKnownFlagsPReg_8_6; // @[AxiLoadQueue.scala 246:86:@38585.8]
  assign _T_93040 = _T_93039 | storeAddrNotKnownFlagsPReg_8_7; // @[AxiLoadQueue.scala 246:86:@38586.8]
  assign _T_93041 = _T_93040 | storeAddrNotKnownFlagsPReg_8_8; // @[AxiLoadQueue.scala 246:86:@38587.8]
  assign _T_93042 = _T_93041 | storeAddrNotKnownFlagsPReg_8_9; // @[AxiLoadQueue.scala 246:86:@38588.8]
  assign _T_93043 = _T_93042 | storeAddrNotKnownFlagsPReg_8_10; // @[AxiLoadQueue.scala 246:86:@38589.8]
  assign _T_93044 = _T_93043 | storeAddrNotKnownFlagsPReg_8_11; // @[AxiLoadQueue.scala 246:86:@38590.8]
  assign _T_93045 = _T_93044 | storeAddrNotKnownFlagsPReg_8_12; // @[AxiLoadQueue.scala 246:86:@38591.8]
  assign _T_93046 = _T_93045 | storeAddrNotKnownFlagsPReg_8_13; // @[AxiLoadQueue.scala 246:86:@38592.8]
  assign _T_93047 = _T_93046 | storeAddrNotKnownFlagsPReg_8_14; // @[AxiLoadQueue.scala 246:86:@38593.8]
  assign _T_93048 = _T_93047 | storeAddrNotKnownFlagsPReg_8_15; // @[AxiLoadQueue.scala 246:86:@38594.8]
  assign _T_93050 = _T_93048 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38595.8]
  assign _T_93069 = _T_89392 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38612.8]
  assign _T_93070 = _T_93050 & _T_93069; // @[AxiLoadQueue.scala 246:103:@38613.8]
  assign _GEN_2032 = _T_93031 ? _T_93070 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38578.6]
  assign loadRequest_8 = _T_93023 ? _GEN_2032 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38572.4]
  assign _T_90469 = loadRequest_8 ? 16'h100 : _T_90468; // @[Mux.scala 31:69:@36522.4]
  assign _T_92938 = dataKnownPReg_7 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38488.4]
  assign _T_92939 = addrKnownPReg_7 & _T_92938; // @[AxiLoadQueue.scala 242:38:@38489.4]
  assign _T_92941 = bypassInitiated_7 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38491.6]
  assign _T_92943 = loadInitiated_7 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38492.6]
  assign _T_92944 = _T_92941 & _T_92943; // @[AxiLoadQueue.scala 243:43:@38493.6]
  assign _T_92946 = dataKnown_7 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38494.6]
  assign _T_92947 = _T_92944 & _T_92946; // @[AxiLoadQueue.scala 243:75:@38495.6]
  assign _T_92950 = storeAddrNotKnownFlagsPReg_7_0 | storeAddrNotKnownFlagsPReg_7_1; // @[AxiLoadQueue.scala 246:86:@38498.8]
  assign _T_92951 = _T_92950 | storeAddrNotKnownFlagsPReg_7_2; // @[AxiLoadQueue.scala 246:86:@38499.8]
  assign _T_92952 = _T_92951 | storeAddrNotKnownFlagsPReg_7_3; // @[AxiLoadQueue.scala 246:86:@38500.8]
  assign _T_92953 = _T_92952 | storeAddrNotKnownFlagsPReg_7_4; // @[AxiLoadQueue.scala 246:86:@38501.8]
  assign _T_92954 = _T_92953 | storeAddrNotKnownFlagsPReg_7_5; // @[AxiLoadQueue.scala 246:86:@38502.8]
  assign _T_92955 = _T_92954 | storeAddrNotKnownFlagsPReg_7_6; // @[AxiLoadQueue.scala 246:86:@38503.8]
  assign _T_92956 = _T_92955 | storeAddrNotKnownFlagsPReg_7_7; // @[AxiLoadQueue.scala 246:86:@38504.8]
  assign _T_92957 = _T_92956 | storeAddrNotKnownFlagsPReg_7_8; // @[AxiLoadQueue.scala 246:86:@38505.8]
  assign _T_92958 = _T_92957 | storeAddrNotKnownFlagsPReg_7_9; // @[AxiLoadQueue.scala 246:86:@38506.8]
  assign _T_92959 = _T_92958 | storeAddrNotKnownFlagsPReg_7_10; // @[AxiLoadQueue.scala 246:86:@38507.8]
  assign _T_92960 = _T_92959 | storeAddrNotKnownFlagsPReg_7_11; // @[AxiLoadQueue.scala 246:86:@38508.8]
  assign _T_92961 = _T_92960 | storeAddrNotKnownFlagsPReg_7_12; // @[AxiLoadQueue.scala 246:86:@38509.8]
  assign _T_92962 = _T_92961 | storeAddrNotKnownFlagsPReg_7_13; // @[AxiLoadQueue.scala 246:86:@38510.8]
  assign _T_92963 = _T_92962 | storeAddrNotKnownFlagsPReg_7_14; // @[AxiLoadQueue.scala 246:86:@38511.8]
  assign _T_92964 = _T_92963 | storeAddrNotKnownFlagsPReg_7_15; // @[AxiLoadQueue.scala 246:86:@38512.8]
  assign _T_92966 = _T_92964 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38513.8]
  assign _T_92985 = _T_89256 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38530.8]
  assign _T_92986 = _T_92966 & _T_92985; // @[AxiLoadQueue.scala 246:103:@38531.8]
  assign _GEN_2028 = _T_92947 ? _T_92986 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38496.6]
  assign loadRequest_7 = _T_92939 ? _GEN_2028 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38490.4]
  assign _T_90470 = loadRequest_7 ? 16'h80 : _T_90469; // @[Mux.scala 31:69:@36523.4]
  assign _T_92854 = dataKnownPReg_6 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38406.4]
  assign _T_92855 = addrKnownPReg_6 & _T_92854; // @[AxiLoadQueue.scala 242:38:@38407.4]
  assign _T_92857 = bypassInitiated_6 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38409.6]
  assign _T_92859 = loadInitiated_6 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38410.6]
  assign _T_92860 = _T_92857 & _T_92859; // @[AxiLoadQueue.scala 243:43:@38411.6]
  assign _T_92862 = dataKnown_6 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38412.6]
  assign _T_92863 = _T_92860 & _T_92862; // @[AxiLoadQueue.scala 243:75:@38413.6]
  assign _T_92866 = storeAddrNotKnownFlagsPReg_6_0 | storeAddrNotKnownFlagsPReg_6_1; // @[AxiLoadQueue.scala 246:86:@38416.8]
  assign _T_92867 = _T_92866 | storeAddrNotKnownFlagsPReg_6_2; // @[AxiLoadQueue.scala 246:86:@38417.8]
  assign _T_92868 = _T_92867 | storeAddrNotKnownFlagsPReg_6_3; // @[AxiLoadQueue.scala 246:86:@38418.8]
  assign _T_92869 = _T_92868 | storeAddrNotKnownFlagsPReg_6_4; // @[AxiLoadQueue.scala 246:86:@38419.8]
  assign _T_92870 = _T_92869 | storeAddrNotKnownFlagsPReg_6_5; // @[AxiLoadQueue.scala 246:86:@38420.8]
  assign _T_92871 = _T_92870 | storeAddrNotKnownFlagsPReg_6_6; // @[AxiLoadQueue.scala 246:86:@38421.8]
  assign _T_92872 = _T_92871 | storeAddrNotKnownFlagsPReg_6_7; // @[AxiLoadQueue.scala 246:86:@38422.8]
  assign _T_92873 = _T_92872 | storeAddrNotKnownFlagsPReg_6_8; // @[AxiLoadQueue.scala 246:86:@38423.8]
  assign _T_92874 = _T_92873 | storeAddrNotKnownFlagsPReg_6_9; // @[AxiLoadQueue.scala 246:86:@38424.8]
  assign _T_92875 = _T_92874 | storeAddrNotKnownFlagsPReg_6_10; // @[AxiLoadQueue.scala 246:86:@38425.8]
  assign _T_92876 = _T_92875 | storeAddrNotKnownFlagsPReg_6_11; // @[AxiLoadQueue.scala 246:86:@38426.8]
  assign _T_92877 = _T_92876 | storeAddrNotKnownFlagsPReg_6_12; // @[AxiLoadQueue.scala 246:86:@38427.8]
  assign _T_92878 = _T_92877 | storeAddrNotKnownFlagsPReg_6_13; // @[AxiLoadQueue.scala 246:86:@38428.8]
  assign _T_92879 = _T_92878 | storeAddrNotKnownFlagsPReg_6_14; // @[AxiLoadQueue.scala 246:86:@38429.8]
  assign _T_92880 = _T_92879 | storeAddrNotKnownFlagsPReg_6_15; // @[AxiLoadQueue.scala 246:86:@38430.8]
  assign _T_92882 = _T_92880 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38431.8]
  assign _T_92901 = _T_89120 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38448.8]
  assign _T_92902 = _T_92882 & _T_92901; // @[AxiLoadQueue.scala 246:103:@38449.8]
  assign _GEN_2024 = _T_92863 ? _T_92902 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38414.6]
  assign loadRequest_6 = _T_92855 ? _GEN_2024 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38408.4]
  assign _T_90471 = loadRequest_6 ? 16'h40 : _T_90470; // @[Mux.scala 31:69:@36524.4]
  assign _T_92770 = dataKnownPReg_5 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38324.4]
  assign _T_92771 = addrKnownPReg_5 & _T_92770; // @[AxiLoadQueue.scala 242:38:@38325.4]
  assign _T_92773 = bypassInitiated_5 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38327.6]
  assign _T_92775 = loadInitiated_5 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38328.6]
  assign _T_92776 = _T_92773 & _T_92775; // @[AxiLoadQueue.scala 243:43:@38329.6]
  assign _T_92778 = dataKnown_5 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38330.6]
  assign _T_92779 = _T_92776 & _T_92778; // @[AxiLoadQueue.scala 243:75:@38331.6]
  assign _T_92782 = storeAddrNotKnownFlagsPReg_5_0 | storeAddrNotKnownFlagsPReg_5_1; // @[AxiLoadQueue.scala 246:86:@38334.8]
  assign _T_92783 = _T_92782 | storeAddrNotKnownFlagsPReg_5_2; // @[AxiLoadQueue.scala 246:86:@38335.8]
  assign _T_92784 = _T_92783 | storeAddrNotKnownFlagsPReg_5_3; // @[AxiLoadQueue.scala 246:86:@38336.8]
  assign _T_92785 = _T_92784 | storeAddrNotKnownFlagsPReg_5_4; // @[AxiLoadQueue.scala 246:86:@38337.8]
  assign _T_92786 = _T_92785 | storeAddrNotKnownFlagsPReg_5_5; // @[AxiLoadQueue.scala 246:86:@38338.8]
  assign _T_92787 = _T_92786 | storeAddrNotKnownFlagsPReg_5_6; // @[AxiLoadQueue.scala 246:86:@38339.8]
  assign _T_92788 = _T_92787 | storeAddrNotKnownFlagsPReg_5_7; // @[AxiLoadQueue.scala 246:86:@38340.8]
  assign _T_92789 = _T_92788 | storeAddrNotKnownFlagsPReg_5_8; // @[AxiLoadQueue.scala 246:86:@38341.8]
  assign _T_92790 = _T_92789 | storeAddrNotKnownFlagsPReg_5_9; // @[AxiLoadQueue.scala 246:86:@38342.8]
  assign _T_92791 = _T_92790 | storeAddrNotKnownFlagsPReg_5_10; // @[AxiLoadQueue.scala 246:86:@38343.8]
  assign _T_92792 = _T_92791 | storeAddrNotKnownFlagsPReg_5_11; // @[AxiLoadQueue.scala 246:86:@38344.8]
  assign _T_92793 = _T_92792 | storeAddrNotKnownFlagsPReg_5_12; // @[AxiLoadQueue.scala 246:86:@38345.8]
  assign _T_92794 = _T_92793 | storeAddrNotKnownFlagsPReg_5_13; // @[AxiLoadQueue.scala 246:86:@38346.8]
  assign _T_92795 = _T_92794 | storeAddrNotKnownFlagsPReg_5_14; // @[AxiLoadQueue.scala 246:86:@38347.8]
  assign _T_92796 = _T_92795 | storeAddrNotKnownFlagsPReg_5_15; // @[AxiLoadQueue.scala 246:86:@38348.8]
  assign _T_92798 = _T_92796 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38349.8]
  assign _T_92817 = _T_88984 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38366.8]
  assign _T_92818 = _T_92798 & _T_92817; // @[AxiLoadQueue.scala 246:103:@38367.8]
  assign _GEN_2020 = _T_92779 ? _T_92818 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38332.6]
  assign loadRequest_5 = _T_92771 ? _GEN_2020 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38326.4]
  assign _T_90472 = loadRequest_5 ? 16'h20 : _T_90471; // @[Mux.scala 31:69:@36525.4]
  assign _T_92686 = dataKnownPReg_4 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38242.4]
  assign _T_92687 = addrKnownPReg_4 & _T_92686; // @[AxiLoadQueue.scala 242:38:@38243.4]
  assign _T_92689 = bypassInitiated_4 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38245.6]
  assign _T_92691 = loadInitiated_4 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38246.6]
  assign _T_92692 = _T_92689 & _T_92691; // @[AxiLoadQueue.scala 243:43:@38247.6]
  assign _T_92694 = dataKnown_4 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38248.6]
  assign _T_92695 = _T_92692 & _T_92694; // @[AxiLoadQueue.scala 243:75:@38249.6]
  assign _T_92698 = storeAddrNotKnownFlagsPReg_4_0 | storeAddrNotKnownFlagsPReg_4_1; // @[AxiLoadQueue.scala 246:86:@38252.8]
  assign _T_92699 = _T_92698 | storeAddrNotKnownFlagsPReg_4_2; // @[AxiLoadQueue.scala 246:86:@38253.8]
  assign _T_92700 = _T_92699 | storeAddrNotKnownFlagsPReg_4_3; // @[AxiLoadQueue.scala 246:86:@38254.8]
  assign _T_92701 = _T_92700 | storeAddrNotKnownFlagsPReg_4_4; // @[AxiLoadQueue.scala 246:86:@38255.8]
  assign _T_92702 = _T_92701 | storeAddrNotKnownFlagsPReg_4_5; // @[AxiLoadQueue.scala 246:86:@38256.8]
  assign _T_92703 = _T_92702 | storeAddrNotKnownFlagsPReg_4_6; // @[AxiLoadQueue.scala 246:86:@38257.8]
  assign _T_92704 = _T_92703 | storeAddrNotKnownFlagsPReg_4_7; // @[AxiLoadQueue.scala 246:86:@38258.8]
  assign _T_92705 = _T_92704 | storeAddrNotKnownFlagsPReg_4_8; // @[AxiLoadQueue.scala 246:86:@38259.8]
  assign _T_92706 = _T_92705 | storeAddrNotKnownFlagsPReg_4_9; // @[AxiLoadQueue.scala 246:86:@38260.8]
  assign _T_92707 = _T_92706 | storeAddrNotKnownFlagsPReg_4_10; // @[AxiLoadQueue.scala 246:86:@38261.8]
  assign _T_92708 = _T_92707 | storeAddrNotKnownFlagsPReg_4_11; // @[AxiLoadQueue.scala 246:86:@38262.8]
  assign _T_92709 = _T_92708 | storeAddrNotKnownFlagsPReg_4_12; // @[AxiLoadQueue.scala 246:86:@38263.8]
  assign _T_92710 = _T_92709 | storeAddrNotKnownFlagsPReg_4_13; // @[AxiLoadQueue.scala 246:86:@38264.8]
  assign _T_92711 = _T_92710 | storeAddrNotKnownFlagsPReg_4_14; // @[AxiLoadQueue.scala 246:86:@38265.8]
  assign _T_92712 = _T_92711 | storeAddrNotKnownFlagsPReg_4_15; // @[AxiLoadQueue.scala 246:86:@38266.8]
  assign _T_92714 = _T_92712 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38267.8]
  assign _T_92733 = _T_88848 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38284.8]
  assign _T_92734 = _T_92714 & _T_92733; // @[AxiLoadQueue.scala 246:103:@38285.8]
  assign _GEN_2016 = _T_92695 ? _T_92734 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38250.6]
  assign loadRequest_4 = _T_92687 ? _GEN_2016 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38244.4]
  assign _T_90473 = loadRequest_4 ? 16'h10 : _T_90472; // @[Mux.scala 31:69:@36526.4]
  assign _T_92602 = dataKnownPReg_3 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38160.4]
  assign _T_92603 = addrKnownPReg_3 & _T_92602; // @[AxiLoadQueue.scala 242:38:@38161.4]
  assign _T_92605 = bypassInitiated_3 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38163.6]
  assign _T_92607 = loadInitiated_3 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38164.6]
  assign _T_92608 = _T_92605 & _T_92607; // @[AxiLoadQueue.scala 243:43:@38165.6]
  assign _T_92610 = dataKnown_3 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38166.6]
  assign _T_92611 = _T_92608 & _T_92610; // @[AxiLoadQueue.scala 243:75:@38167.6]
  assign _T_92614 = storeAddrNotKnownFlagsPReg_3_0 | storeAddrNotKnownFlagsPReg_3_1; // @[AxiLoadQueue.scala 246:86:@38170.8]
  assign _T_92615 = _T_92614 | storeAddrNotKnownFlagsPReg_3_2; // @[AxiLoadQueue.scala 246:86:@38171.8]
  assign _T_92616 = _T_92615 | storeAddrNotKnownFlagsPReg_3_3; // @[AxiLoadQueue.scala 246:86:@38172.8]
  assign _T_92617 = _T_92616 | storeAddrNotKnownFlagsPReg_3_4; // @[AxiLoadQueue.scala 246:86:@38173.8]
  assign _T_92618 = _T_92617 | storeAddrNotKnownFlagsPReg_3_5; // @[AxiLoadQueue.scala 246:86:@38174.8]
  assign _T_92619 = _T_92618 | storeAddrNotKnownFlagsPReg_3_6; // @[AxiLoadQueue.scala 246:86:@38175.8]
  assign _T_92620 = _T_92619 | storeAddrNotKnownFlagsPReg_3_7; // @[AxiLoadQueue.scala 246:86:@38176.8]
  assign _T_92621 = _T_92620 | storeAddrNotKnownFlagsPReg_3_8; // @[AxiLoadQueue.scala 246:86:@38177.8]
  assign _T_92622 = _T_92621 | storeAddrNotKnownFlagsPReg_3_9; // @[AxiLoadQueue.scala 246:86:@38178.8]
  assign _T_92623 = _T_92622 | storeAddrNotKnownFlagsPReg_3_10; // @[AxiLoadQueue.scala 246:86:@38179.8]
  assign _T_92624 = _T_92623 | storeAddrNotKnownFlagsPReg_3_11; // @[AxiLoadQueue.scala 246:86:@38180.8]
  assign _T_92625 = _T_92624 | storeAddrNotKnownFlagsPReg_3_12; // @[AxiLoadQueue.scala 246:86:@38181.8]
  assign _T_92626 = _T_92625 | storeAddrNotKnownFlagsPReg_3_13; // @[AxiLoadQueue.scala 246:86:@38182.8]
  assign _T_92627 = _T_92626 | storeAddrNotKnownFlagsPReg_3_14; // @[AxiLoadQueue.scala 246:86:@38183.8]
  assign _T_92628 = _T_92627 | storeAddrNotKnownFlagsPReg_3_15; // @[AxiLoadQueue.scala 246:86:@38184.8]
  assign _T_92630 = _T_92628 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38185.8]
  assign _T_92649 = _T_88712 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38202.8]
  assign _T_92650 = _T_92630 & _T_92649; // @[AxiLoadQueue.scala 246:103:@38203.8]
  assign _GEN_2012 = _T_92611 ? _T_92650 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38168.6]
  assign loadRequest_3 = _T_92603 ? _GEN_2012 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38162.4]
  assign _T_90474 = loadRequest_3 ? 16'h8 : _T_90473; // @[Mux.scala 31:69:@36527.4]
  assign _T_92518 = dataKnownPReg_2 == 1'h0; // @[AxiLoadQueue.scala 242:41:@38078.4]
  assign _T_92519 = addrKnownPReg_2 & _T_92518; // @[AxiLoadQueue.scala 242:38:@38079.4]
  assign _T_92521 = bypassInitiated_2 == 1'h0; // @[AxiLoadQueue.scala 243:12:@38081.6]
  assign _T_92523 = loadInitiated_2 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38082.6]
  assign _T_92524 = _T_92521 & _T_92523; // @[AxiLoadQueue.scala 243:43:@38083.6]
  assign _T_92526 = dataKnown_2 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38084.6]
  assign _T_92527 = _T_92524 & _T_92526; // @[AxiLoadQueue.scala 243:75:@38085.6]
  assign _T_92530 = storeAddrNotKnownFlagsPReg_2_0 | storeAddrNotKnownFlagsPReg_2_1; // @[AxiLoadQueue.scala 246:86:@38088.8]
  assign _T_92531 = _T_92530 | storeAddrNotKnownFlagsPReg_2_2; // @[AxiLoadQueue.scala 246:86:@38089.8]
  assign _T_92532 = _T_92531 | storeAddrNotKnownFlagsPReg_2_3; // @[AxiLoadQueue.scala 246:86:@38090.8]
  assign _T_92533 = _T_92532 | storeAddrNotKnownFlagsPReg_2_4; // @[AxiLoadQueue.scala 246:86:@38091.8]
  assign _T_92534 = _T_92533 | storeAddrNotKnownFlagsPReg_2_5; // @[AxiLoadQueue.scala 246:86:@38092.8]
  assign _T_92535 = _T_92534 | storeAddrNotKnownFlagsPReg_2_6; // @[AxiLoadQueue.scala 246:86:@38093.8]
  assign _T_92536 = _T_92535 | storeAddrNotKnownFlagsPReg_2_7; // @[AxiLoadQueue.scala 246:86:@38094.8]
  assign _T_92537 = _T_92536 | storeAddrNotKnownFlagsPReg_2_8; // @[AxiLoadQueue.scala 246:86:@38095.8]
  assign _T_92538 = _T_92537 | storeAddrNotKnownFlagsPReg_2_9; // @[AxiLoadQueue.scala 246:86:@38096.8]
  assign _T_92539 = _T_92538 | storeAddrNotKnownFlagsPReg_2_10; // @[AxiLoadQueue.scala 246:86:@38097.8]
  assign _T_92540 = _T_92539 | storeAddrNotKnownFlagsPReg_2_11; // @[AxiLoadQueue.scala 246:86:@38098.8]
  assign _T_92541 = _T_92540 | storeAddrNotKnownFlagsPReg_2_12; // @[AxiLoadQueue.scala 246:86:@38099.8]
  assign _T_92542 = _T_92541 | storeAddrNotKnownFlagsPReg_2_13; // @[AxiLoadQueue.scala 246:86:@38100.8]
  assign _T_92543 = _T_92542 | storeAddrNotKnownFlagsPReg_2_14; // @[AxiLoadQueue.scala 246:86:@38101.8]
  assign _T_92544 = _T_92543 | storeAddrNotKnownFlagsPReg_2_15; // @[AxiLoadQueue.scala 246:86:@38102.8]
  assign _T_92546 = _T_92544 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38103.8]
  assign _T_92565 = _T_88576 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38120.8]
  assign _T_92566 = _T_92546 & _T_92565; // @[AxiLoadQueue.scala 246:103:@38121.8]
  assign _GEN_2008 = _T_92527 ? _T_92566 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38086.6]
  assign loadRequest_2 = _T_92519 ? _GEN_2008 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38080.4]
  assign _T_90475 = loadRequest_2 ? 16'h4 : _T_90474; // @[Mux.scala 31:69:@36528.4]
  assign _T_92434 = dataKnownPReg_1 == 1'h0; // @[AxiLoadQueue.scala 242:41:@37996.4]
  assign _T_92435 = addrKnownPReg_1 & _T_92434; // @[AxiLoadQueue.scala 242:38:@37997.4]
  assign _T_92437 = bypassInitiated_1 == 1'h0; // @[AxiLoadQueue.scala 243:12:@37999.6]
  assign _T_92439 = loadInitiated_1 == 1'h0; // @[AxiLoadQueue.scala 243:46:@38000.6]
  assign _T_92440 = _T_92437 & _T_92439; // @[AxiLoadQueue.scala 243:43:@38001.6]
  assign _T_92442 = dataKnown_1 == 1'h0; // @[AxiLoadQueue.scala 243:78:@38002.6]
  assign _T_92443 = _T_92440 & _T_92442; // @[AxiLoadQueue.scala 243:75:@38003.6]
  assign _T_92446 = storeAddrNotKnownFlagsPReg_1_0 | storeAddrNotKnownFlagsPReg_1_1; // @[AxiLoadQueue.scala 246:86:@38006.8]
  assign _T_92447 = _T_92446 | storeAddrNotKnownFlagsPReg_1_2; // @[AxiLoadQueue.scala 246:86:@38007.8]
  assign _T_92448 = _T_92447 | storeAddrNotKnownFlagsPReg_1_3; // @[AxiLoadQueue.scala 246:86:@38008.8]
  assign _T_92449 = _T_92448 | storeAddrNotKnownFlagsPReg_1_4; // @[AxiLoadQueue.scala 246:86:@38009.8]
  assign _T_92450 = _T_92449 | storeAddrNotKnownFlagsPReg_1_5; // @[AxiLoadQueue.scala 246:86:@38010.8]
  assign _T_92451 = _T_92450 | storeAddrNotKnownFlagsPReg_1_6; // @[AxiLoadQueue.scala 246:86:@38011.8]
  assign _T_92452 = _T_92451 | storeAddrNotKnownFlagsPReg_1_7; // @[AxiLoadQueue.scala 246:86:@38012.8]
  assign _T_92453 = _T_92452 | storeAddrNotKnownFlagsPReg_1_8; // @[AxiLoadQueue.scala 246:86:@38013.8]
  assign _T_92454 = _T_92453 | storeAddrNotKnownFlagsPReg_1_9; // @[AxiLoadQueue.scala 246:86:@38014.8]
  assign _T_92455 = _T_92454 | storeAddrNotKnownFlagsPReg_1_10; // @[AxiLoadQueue.scala 246:86:@38015.8]
  assign _T_92456 = _T_92455 | storeAddrNotKnownFlagsPReg_1_11; // @[AxiLoadQueue.scala 246:86:@38016.8]
  assign _T_92457 = _T_92456 | storeAddrNotKnownFlagsPReg_1_12; // @[AxiLoadQueue.scala 246:86:@38017.8]
  assign _T_92458 = _T_92457 | storeAddrNotKnownFlagsPReg_1_13; // @[AxiLoadQueue.scala 246:86:@38018.8]
  assign _T_92459 = _T_92458 | storeAddrNotKnownFlagsPReg_1_14; // @[AxiLoadQueue.scala 246:86:@38019.8]
  assign _T_92460 = _T_92459 | storeAddrNotKnownFlagsPReg_1_15; // @[AxiLoadQueue.scala 246:86:@38020.8]
  assign _T_92462 = _T_92460 == 1'h0; // @[AxiLoadQueue.scala 246:38:@38021.8]
  assign _T_92481 = _T_88440 == 1'h0; // @[AxiLoadQueue.scala 247:11:@38038.8]
  assign _T_92482 = _T_92462 & _T_92481; // @[AxiLoadQueue.scala 246:103:@38039.8]
  assign _GEN_2004 = _T_92443 ? _T_92482 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38004.6]
  assign loadRequest_1 = _T_92435 ? _GEN_2004 : 1'h0; // @[AxiLoadQueue.scala 242:71:@37998.4]
  assign _T_90476 = loadRequest_1 ? 16'h2 : _T_90475; // @[Mux.scala 31:69:@36529.4]
  assign _T_92350 = dataKnownPReg_0 == 1'h0; // @[AxiLoadQueue.scala 242:41:@37914.4]
  assign _T_92351 = addrKnownPReg_0 & _T_92350; // @[AxiLoadQueue.scala 242:38:@37915.4]
  assign _T_92353 = bypassInitiated_0 == 1'h0; // @[AxiLoadQueue.scala 243:12:@37917.6]
  assign _T_92355 = loadInitiated_0 == 1'h0; // @[AxiLoadQueue.scala 243:46:@37918.6]
  assign _T_92356 = _T_92353 & _T_92355; // @[AxiLoadQueue.scala 243:43:@37919.6]
  assign _T_92358 = dataKnown_0 == 1'h0; // @[AxiLoadQueue.scala 243:78:@37920.6]
  assign _T_92359 = _T_92356 & _T_92358; // @[AxiLoadQueue.scala 243:75:@37921.6]
  assign _T_92362 = storeAddrNotKnownFlagsPReg_0_0 | storeAddrNotKnownFlagsPReg_0_1; // @[AxiLoadQueue.scala 246:86:@37924.8]
  assign _T_92363 = _T_92362 | storeAddrNotKnownFlagsPReg_0_2; // @[AxiLoadQueue.scala 246:86:@37925.8]
  assign _T_92364 = _T_92363 | storeAddrNotKnownFlagsPReg_0_3; // @[AxiLoadQueue.scala 246:86:@37926.8]
  assign _T_92365 = _T_92364 | storeAddrNotKnownFlagsPReg_0_4; // @[AxiLoadQueue.scala 246:86:@37927.8]
  assign _T_92366 = _T_92365 | storeAddrNotKnownFlagsPReg_0_5; // @[AxiLoadQueue.scala 246:86:@37928.8]
  assign _T_92367 = _T_92366 | storeAddrNotKnownFlagsPReg_0_6; // @[AxiLoadQueue.scala 246:86:@37929.8]
  assign _T_92368 = _T_92367 | storeAddrNotKnownFlagsPReg_0_7; // @[AxiLoadQueue.scala 246:86:@37930.8]
  assign _T_92369 = _T_92368 | storeAddrNotKnownFlagsPReg_0_8; // @[AxiLoadQueue.scala 246:86:@37931.8]
  assign _T_92370 = _T_92369 | storeAddrNotKnownFlagsPReg_0_9; // @[AxiLoadQueue.scala 246:86:@37932.8]
  assign _T_92371 = _T_92370 | storeAddrNotKnownFlagsPReg_0_10; // @[AxiLoadQueue.scala 246:86:@37933.8]
  assign _T_92372 = _T_92371 | storeAddrNotKnownFlagsPReg_0_11; // @[AxiLoadQueue.scala 246:86:@37934.8]
  assign _T_92373 = _T_92372 | storeAddrNotKnownFlagsPReg_0_12; // @[AxiLoadQueue.scala 246:86:@37935.8]
  assign _T_92374 = _T_92373 | storeAddrNotKnownFlagsPReg_0_13; // @[AxiLoadQueue.scala 246:86:@37936.8]
  assign _T_92375 = _T_92374 | storeAddrNotKnownFlagsPReg_0_14; // @[AxiLoadQueue.scala 246:86:@37937.8]
  assign _T_92376 = _T_92375 | storeAddrNotKnownFlagsPReg_0_15; // @[AxiLoadQueue.scala 246:86:@37938.8]
  assign _T_92378 = _T_92376 == 1'h0; // @[AxiLoadQueue.scala 246:38:@37939.8]
  assign _T_92397 = _T_88304 == 1'h0; // @[AxiLoadQueue.scala 247:11:@37956.8]
  assign _T_92398 = _T_92378 & _T_92397; // @[AxiLoadQueue.scala 246:103:@37957.8]
  assign _GEN_2000 = _T_92359 ? _T_92398 : 1'h0; // @[AxiLoadQueue.scala 243:104:@37922.6]
  assign loadRequest_0 = _T_92351 ? _GEN_2000 : 1'h0; // @[AxiLoadQueue.scala 242:71:@37916.4]
  assign _T_90477 = loadRequest_0 ? 16'h1 : _T_90476; // @[Mux.scala 31:69:@36530.4]
  assign _T_90478 = _T_90477[0]; // @[OneHot.scala 66:30:@36531.4]
  assign _T_90479 = _T_90477[1]; // @[OneHot.scala 66:30:@36532.4]
  assign _T_90480 = _T_90477[2]; // @[OneHot.scala 66:30:@36533.4]
  assign _T_90481 = _T_90477[3]; // @[OneHot.scala 66:30:@36534.4]
  assign _T_90482 = _T_90477[4]; // @[OneHot.scala 66:30:@36535.4]
  assign _T_90483 = _T_90477[5]; // @[OneHot.scala 66:30:@36536.4]
  assign _T_90484 = _T_90477[6]; // @[OneHot.scala 66:30:@36537.4]
  assign _T_90485 = _T_90477[7]; // @[OneHot.scala 66:30:@36538.4]
  assign _T_90486 = _T_90477[8]; // @[OneHot.scala 66:30:@36539.4]
  assign _T_90487 = _T_90477[9]; // @[OneHot.scala 66:30:@36540.4]
  assign _T_90488 = _T_90477[10]; // @[OneHot.scala 66:30:@36541.4]
  assign _T_90489 = _T_90477[11]; // @[OneHot.scala 66:30:@36542.4]
  assign _T_90490 = _T_90477[12]; // @[OneHot.scala 66:30:@36543.4]
  assign _T_90491 = _T_90477[13]; // @[OneHot.scala 66:30:@36544.4]
  assign _T_90492 = _T_90477[14]; // @[OneHot.scala 66:30:@36545.4]
  assign _T_90493 = _T_90477[15]; // @[OneHot.scala 66:30:@36546.4]
  assign _T_90534 = loadRequest_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36564.4]
  assign _T_90535 = loadRequest_15 ? 16'h4000 : _T_90534; // @[Mux.scala 31:69:@36565.4]
  assign _T_90536 = loadRequest_14 ? 16'h2000 : _T_90535; // @[Mux.scala 31:69:@36566.4]
  assign _T_90537 = loadRequest_13 ? 16'h1000 : _T_90536; // @[Mux.scala 31:69:@36567.4]
  assign _T_90538 = loadRequest_12 ? 16'h800 : _T_90537; // @[Mux.scala 31:69:@36568.4]
  assign _T_90539 = loadRequest_11 ? 16'h400 : _T_90538; // @[Mux.scala 31:69:@36569.4]
  assign _T_90540 = loadRequest_10 ? 16'h200 : _T_90539; // @[Mux.scala 31:69:@36570.4]
  assign _T_90541 = loadRequest_9 ? 16'h100 : _T_90540; // @[Mux.scala 31:69:@36571.4]
  assign _T_90542 = loadRequest_8 ? 16'h80 : _T_90541; // @[Mux.scala 31:69:@36572.4]
  assign _T_90543 = loadRequest_7 ? 16'h40 : _T_90542; // @[Mux.scala 31:69:@36573.4]
  assign _T_90544 = loadRequest_6 ? 16'h20 : _T_90543; // @[Mux.scala 31:69:@36574.4]
  assign _T_90545 = loadRequest_5 ? 16'h10 : _T_90544; // @[Mux.scala 31:69:@36575.4]
  assign _T_90546 = loadRequest_4 ? 16'h8 : _T_90545; // @[Mux.scala 31:69:@36576.4]
  assign _T_90547 = loadRequest_3 ? 16'h4 : _T_90546; // @[Mux.scala 31:69:@36577.4]
  assign _T_90548 = loadRequest_2 ? 16'h2 : _T_90547; // @[Mux.scala 31:69:@36578.4]
  assign _T_90549 = loadRequest_1 ? 16'h1 : _T_90548; // @[Mux.scala 31:69:@36579.4]
  assign _T_90550 = _T_90549[0]; // @[OneHot.scala 66:30:@36580.4]
  assign _T_90551 = _T_90549[1]; // @[OneHot.scala 66:30:@36581.4]
  assign _T_90552 = _T_90549[2]; // @[OneHot.scala 66:30:@36582.4]
  assign _T_90553 = _T_90549[3]; // @[OneHot.scala 66:30:@36583.4]
  assign _T_90554 = _T_90549[4]; // @[OneHot.scala 66:30:@36584.4]
  assign _T_90555 = _T_90549[5]; // @[OneHot.scala 66:30:@36585.4]
  assign _T_90556 = _T_90549[6]; // @[OneHot.scala 66:30:@36586.4]
  assign _T_90557 = _T_90549[7]; // @[OneHot.scala 66:30:@36587.4]
  assign _T_90558 = _T_90549[8]; // @[OneHot.scala 66:30:@36588.4]
  assign _T_90559 = _T_90549[9]; // @[OneHot.scala 66:30:@36589.4]
  assign _T_90560 = _T_90549[10]; // @[OneHot.scala 66:30:@36590.4]
  assign _T_90561 = _T_90549[11]; // @[OneHot.scala 66:30:@36591.4]
  assign _T_90562 = _T_90549[12]; // @[OneHot.scala 66:30:@36592.4]
  assign _T_90563 = _T_90549[13]; // @[OneHot.scala 66:30:@36593.4]
  assign _T_90564 = _T_90549[14]; // @[OneHot.scala 66:30:@36594.4]
  assign _T_90565 = _T_90549[15]; // @[OneHot.scala 66:30:@36595.4]
  assign _T_90606 = loadRequest_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36613.4]
  assign _T_90607 = loadRequest_0 ? 16'h4000 : _T_90606; // @[Mux.scala 31:69:@36614.4]
  assign _T_90608 = loadRequest_15 ? 16'h2000 : _T_90607; // @[Mux.scala 31:69:@36615.4]
  assign _T_90609 = loadRequest_14 ? 16'h1000 : _T_90608; // @[Mux.scala 31:69:@36616.4]
  assign _T_90610 = loadRequest_13 ? 16'h800 : _T_90609; // @[Mux.scala 31:69:@36617.4]
  assign _T_90611 = loadRequest_12 ? 16'h400 : _T_90610; // @[Mux.scala 31:69:@36618.4]
  assign _T_90612 = loadRequest_11 ? 16'h200 : _T_90611; // @[Mux.scala 31:69:@36619.4]
  assign _T_90613 = loadRequest_10 ? 16'h100 : _T_90612; // @[Mux.scala 31:69:@36620.4]
  assign _T_90614 = loadRequest_9 ? 16'h80 : _T_90613; // @[Mux.scala 31:69:@36621.4]
  assign _T_90615 = loadRequest_8 ? 16'h40 : _T_90614; // @[Mux.scala 31:69:@36622.4]
  assign _T_90616 = loadRequest_7 ? 16'h20 : _T_90615; // @[Mux.scala 31:69:@36623.4]
  assign _T_90617 = loadRequest_6 ? 16'h10 : _T_90616; // @[Mux.scala 31:69:@36624.4]
  assign _T_90618 = loadRequest_5 ? 16'h8 : _T_90617; // @[Mux.scala 31:69:@36625.4]
  assign _T_90619 = loadRequest_4 ? 16'h4 : _T_90618; // @[Mux.scala 31:69:@36626.4]
  assign _T_90620 = loadRequest_3 ? 16'h2 : _T_90619; // @[Mux.scala 31:69:@36627.4]
  assign _T_90621 = loadRequest_2 ? 16'h1 : _T_90620; // @[Mux.scala 31:69:@36628.4]
  assign _T_90622 = _T_90621[0]; // @[OneHot.scala 66:30:@36629.4]
  assign _T_90623 = _T_90621[1]; // @[OneHot.scala 66:30:@36630.4]
  assign _T_90624 = _T_90621[2]; // @[OneHot.scala 66:30:@36631.4]
  assign _T_90625 = _T_90621[3]; // @[OneHot.scala 66:30:@36632.4]
  assign _T_90626 = _T_90621[4]; // @[OneHot.scala 66:30:@36633.4]
  assign _T_90627 = _T_90621[5]; // @[OneHot.scala 66:30:@36634.4]
  assign _T_90628 = _T_90621[6]; // @[OneHot.scala 66:30:@36635.4]
  assign _T_90629 = _T_90621[7]; // @[OneHot.scala 66:30:@36636.4]
  assign _T_90630 = _T_90621[8]; // @[OneHot.scala 66:30:@36637.4]
  assign _T_90631 = _T_90621[9]; // @[OneHot.scala 66:30:@36638.4]
  assign _T_90632 = _T_90621[10]; // @[OneHot.scala 66:30:@36639.4]
  assign _T_90633 = _T_90621[11]; // @[OneHot.scala 66:30:@36640.4]
  assign _T_90634 = _T_90621[12]; // @[OneHot.scala 66:30:@36641.4]
  assign _T_90635 = _T_90621[13]; // @[OneHot.scala 66:30:@36642.4]
  assign _T_90636 = _T_90621[14]; // @[OneHot.scala 66:30:@36643.4]
  assign _T_90637 = _T_90621[15]; // @[OneHot.scala 66:30:@36644.4]
  assign _T_90678 = loadRequest_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36662.4]
  assign _T_90679 = loadRequest_1 ? 16'h4000 : _T_90678; // @[Mux.scala 31:69:@36663.4]
  assign _T_90680 = loadRequest_0 ? 16'h2000 : _T_90679; // @[Mux.scala 31:69:@36664.4]
  assign _T_90681 = loadRequest_15 ? 16'h1000 : _T_90680; // @[Mux.scala 31:69:@36665.4]
  assign _T_90682 = loadRequest_14 ? 16'h800 : _T_90681; // @[Mux.scala 31:69:@36666.4]
  assign _T_90683 = loadRequest_13 ? 16'h400 : _T_90682; // @[Mux.scala 31:69:@36667.4]
  assign _T_90684 = loadRequest_12 ? 16'h200 : _T_90683; // @[Mux.scala 31:69:@36668.4]
  assign _T_90685 = loadRequest_11 ? 16'h100 : _T_90684; // @[Mux.scala 31:69:@36669.4]
  assign _T_90686 = loadRequest_10 ? 16'h80 : _T_90685; // @[Mux.scala 31:69:@36670.4]
  assign _T_90687 = loadRequest_9 ? 16'h40 : _T_90686; // @[Mux.scala 31:69:@36671.4]
  assign _T_90688 = loadRequest_8 ? 16'h20 : _T_90687; // @[Mux.scala 31:69:@36672.4]
  assign _T_90689 = loadRequest_7 ? 16'h10 : _T_90688; // @[Mux.scala 31:69:@36673.4]
  assign _T_90690 = loadRequest_6 ? 16'h8 : _T_90689; // @[Mux.scala 31:69:@36674.4]
  assign _T_90691 = loadRequest_5 ? 16'h4 : _T_90690; // @[Mux.scala 31:69:@36675.4]
  assign _T_90692 = loadRequest_4 ? 16'h2 : _T_90691; // @[Mux.scala 31:69:@36676.4]
  assign _T_90693 = loadRequest_3 ? 16'h1 : _T_90692; // @[Mux.scala 31:69:@36677.4]
  assign _T_90694 = _T_90693[0]; // @[OneHot.scala 66:30:@36678.4]
  assign _T_90695 = _T_90693[1]; // @[OneHot.scala 66:30:@36679.4]
  assign _T_90696 = _T_90693[2]; // @[OneHot.scala 66:30:@36680.4]
  assign _T_90697 = _T_90693[3]; // @[OneHot.scala 66:30:@36681.4]
  assign _T_90698 = _T_90693[4]; // @[OneHot.scala 66:30:@36682.4]
  assign _T_90699 = _T_90693[5]; // @[OneHot.scala 66:30:@36683.4]
  assign _T_90700 = _T_90693[6]; // @[OneHot.scala 66:30:@36684.4]
  assign _T_90701 = _T_90693[7]; // @[OneHot.scala 66:30:@36685.4]
  assign _T_90702 = _T_90693[8]; // @[OneHot.scala 66:30:@36686.4]
  assign _T_90703 = _T_90693[9]; // @[OneHot.scala 66:30:@36687.4]
  assign _T_90704 = _T_90693[10]; // @[OneHot.scala 66:30:@36688.4]
  assign _T_90705 = _T_90693[11]; // @[OneHot.scala 66:30:@36689.4]
  assign _T_90706 = _T_90693[12]; // @[OneHot.scala 66:30:@36690.4]
  assign _T_90707 = _T_90693[13]; // @[OneHot.scala 66:30:@36691.4]
  assign _T_90708 = _T_90693[14]; // @[OneHot.scala 66:30:@36692.4]
  assign _T_90709 = _T_90693[15]; // @[OneHot.scala 66:30:@36693.4]
  assign _T_90750 = loadRequest_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36711.4]
  assign _T_90751 = loadRequest_2 ? 16'h4000 : _T_90750; // @[Mux.scala 31:69:@36712.4]
  assign _T_90752 = loadRequest_1 ? 16'h2000 : _T_90751; // @[Mux.scala 31:69:@36713.4]
  assign _T_90753 = loadRequest_0 ? 16'h1000 : _T_90752; // @[Mux.scala 31:69:@36714.4]
  assign _T_90754 = loadRequest_15 ? 16'h800 : _T_90753; // @[Mux.scala 31:69:@36715.4]
  assign _T_90755 = loadRequest_14 ? 16'h400 : _T_90754; // @[Mux.scala 31:69:@36716.4]
  assign _T_90756 = loadRequest_13 ? 16'h200 : _T_90755; // @[Mux.scala 31:69:@36717.4]
  assign _T_90757 = loadRequest_12 ? 16'h100 : _T_90756; // @[Mux.scala 31:69:@36718.4]
  assign _T_90758 = loadRequest_11 ? 16'h80 : _T_90757; // @[Mux.scala 31:69:@36719.4]
  assign _T_90759 = loadRequest_10 ? 16'h40 : _T_90758; // @[Mux.scala 31:69:@36720.4]
  assign _T_90760 = loadRequest_9 ? 16'h20 : _T_90759; // @[Mux.scala 31:69:@36721.4]
  assign _T_90761 = loadRequest_8 ? 16'h10 : _T_90760; // @[Mux.scala 31:69:@36722.4]
  assign _T_90762 = loadRequest_7 ? 16'h8 : _T_90761; // @[Mux.scala 31:69:@36723.4]
  assign _T_90763 = loadRequest_6 ? 16'h4 : _T_90762; // @[Mux.scala 31:69:@36724.4]
  assign _T_90764 = loadRequest_5 ? 16'h2 : _T_90763; // @[Mux.scala 31:69:@36725.4]
  assign _T_90765 = loadRequest_4 ? 16'h1 : _T_90764; // @[Mux.scala 31:69:@36726.4]
  assign _T_90766 = _T_90765[0]; // @[OneHot.scala 66:30:@36727.4]
  assign _T_90767 = _T_90765[1]; // @[OneHot.scala 66:30:@36728.4]
  assign _T_90768 = _T_90765[2]; // @[OneHot.scala 66:30:@36729.4]
  assign _T_90769 = _T_90765[3]; // @[OneHot.scala 66:30:@36730.4]
  assign _T_90770 = _T_90765[4]; // @[OneHot.scala 66:30:@36731.4]
  assign _T_90771 = _T_90765[5]; // @[OneHot.scala 66:30:@36732.4]
  assign _T_90772 = _T_90765[6]; // @[OneHot.scala 66:30:@36733.4]
  assign _T_90773 = _T_90765[7]; // @[OneHot.scala 66:30:@36734.4]
  assign _T_90774 = _T_90765[8]; // @[OneHot.scala 66:30:@36735.4]
  assign _T_90775 = _T_90765[9]; // @[OneHot.scala 66:30:@36736.4]
  assign _T_90776 = _T_90765[10]; // @[OneHot.scala 66:30:@36737.4]
  assign _T_90777 = _T_90765[11]; // @[OneHot.scala 66:30:@36738.4]
  assign _T_90778 = _T_90765[12]; // @[OneHot.scala 66:30:@36739.4]
  assign _T_90779 = _T_90765[13]; // @[OneHot.scala 66:30:@36740.4]
  assign _T_90780 = _T_90765[14]; // @[OneHot.scala 66:30:@36741.4]
  assign _T_90781 = _T_90765[15]; // @[OneHot.scala 66:30:@36742.4]
  assign _T_90822 = loadRequest_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36760.4]
  assign _T_90823 = loadRequest_3 ? 16'h4000 : _T_90822; // @[Mux.scala 31:69:@36761.4]
  assign _T_90824 = loadRequest_2 ? 16'h2000 : _T_90823; // @[Mux.scala 31:69:@36762.4]
  assign _T_90825 = loadRequest_1 ? 16'h1000 : _T_90824; // @[Mux.scala 31:69:@36763.4]
  assign _T_90826 = loadRequest_0 ? 16'h800 : _T_90825; // @[Mux.scala 31:69:@36764.4]
  assign _T_90827 = loadRequest_15 ? 16'h400 : _T_90826; // @[Mux.scala 31:69:@36765.4]
  assign _T_90828 = loadRequest_14 ? 16'h200 : _T_90827; // @[Mux.scala 31:69:@36766.4]
  assign _T_90829 = loadRequest_13 ? 16'h100 : _T_90828; // @[Mux.scala 31:69:@36767.4]
  assign _T_90830 = loadRequest_12 ? 16'h80 : _T_90829; // @[Mux.scala 31:69:@36768.4]
  assign _T_90831 = loadRequest_11 ? 16'h40 : _T_90830; // @[Mux.scala 31:69:@36769.4]
  assign _T_90832 = loadRequest_10 ? 16'h20 : _T_90831; // @[Mux.scala 31:69:@36770.4]
  assign _T_90833 = loadRequest_9 ? 16'h10 : _T_90832; // @[Mux.scala 31:69:@36771.4]
  assign _T_90834 = loadRequest_8 ? 16'h8 : _T_90833; // @[Mux.scala 31:69:@36772.4]
  assign _T_90835 = loadRequest_7 ? 16'h4 : _T_90834; // @[Mux.scala 31:69:@36773.4]
  assign _T_90836 = loadRequest_6 ? 16'h2 : _T_90835; // @[Mux.scala 31:69:@36774.4]
  assign _T_90837 = loadRequest_5 ? 16'h1 : _T_90836; // @[Mux.scala 31:69:@36775.4]
  assign _T_90838 = _T_90837[0]; // @[OneHot.scala 66:30:@36776.4]
  assign _T_90839 = _T_90837[1]; // @[OneHot.scala 66:30:@36777.4]
  assign _T_90840 = _T_90837[2]; // @[OneHot.scala 66:30:@36778.4]
  assign _T_90841 = _T_90837[3]; // @[OneHot.scala 66:30:@36779.4]
  assign _T_90842 = _T_90837[4]; // @[OneHot.scala 66:30:@36780.4]
  assign _T_90843 = _T_90837[5]; // @[OneHot.scala 66:30:@36781.4]
  assign _T_90844 = _T_90837[6]; // @[OneHot.scala 66:30:@36782.4]
  assign _T_90845 = _T_90837[7]; // @[OneHot.scala 66:30:@36783.4]
  assign _T_90846 = _T_90837[8]; // @[OneHot.scala 66:30:@36784.4]
  assign _T_90847 = _T_90837[9]; // @[OneHot.scala 66:30:@36785.4]
  assign _T_90848 = _T_90837[10]; // @[OneHot.scala 66:30:@36786.4]
  assign _T_90849 = _T_90837[11]; // @[OneHot.scala 66:30:@36787.4]
  assign _T_90850 = _T_90837[12]; // @[OneHot.scala 66:30:@36788.4]
  assign _T_90851 = _T_90837[13]; // @[OneHot.scala 66:30:@36789.4]
  assign _T_90852 = _T_90837[14]; // @[OneHot.scala 66:30:@36790.4]
  assign _T_90853 = _T_90837[15]; // @[OneHot.scala 66:30:@36791.4]
  assign _T_90894 = loadRequest_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36809.4]
  assign _T_90895 = loadRequest_4 ? 16'h4000 : _T_90894; // @[Mux.scala 31:69:@36810.4]
  assign _T_90896 = loadRequest_3 ? 16'h2000 : _T_90895; // @[Mux.scala 31:69:@36811.4]
  assign _T_90897 = loadRequest_2 ? 16'h1000 : _T_90896; // @[Mux.scala 31:69:@36812.4]
  assign _T_90898 = loadRequest_1 ? 16'h800 : _T_90897; // @[Mux.scala 31:69:@36813.4]
  assign _T_90899 = loadRequest_0 ? 16'h400 : _T_90898; // @[Mux.scala 31:69:@36814.4]
  assign _T_90900 = loadRequest_15 ? 16'h200 : _T_90899; // @[Mux.scala 31:69:@36815.4]
  assign _T_90901 = loadRequest_14 ? 16'h100 : _T_90900; // @[Mux.scala 31:69:@36816.4]
  assign _T_90902 = loadRequest_13 ? 16'h80 : _T_90901; // @[Mux.scala 31:69:@36817.4]
  assign _T_90903 = loadRequest_12 ? 16'h40 : _T_90902; // @[Mux.scala 31:69:@36818.4]
  assign _T_90904 = loadRequest_11 ? 16'h20 : _T_90903; // @[Mux.scala 31:69:@36819.4]
  assign _T_90905 = loadRequest_10 ? 16'h10 : _T_90904; // @[Mux.scala 31:69:@36820.4]
  assign _T_90906 = loadRequest_9 ? 16'h8 : _T_90905; // @[Mux.scala 31:69:@36821.4]
  assign _T_90907 = loadRequest_8 ? 16'h4 : _T_90906; // @[Mux.scala 31:69:@36822.4]
  assign _T_90908 = loadRequest_7 ? 16'h2 : _T_90907; // @[Mux.scala 31:69:@36823.4]
  assign _T_90909 = loadRequest_6 ? 16'h1 : _T_90908; // @[Mux.scala 31:69:@36824.4]
  assign _T_90910 = _T_90909[0]; // @[OneHot.scala 66:30:@36825.4]
  assign _T_90911 = _T_90909[1]; // @[OneHot.scala 66:30:@36826.4]
  assign _T_90912 = _T_90909[2]; // @[OneHot.scala 66:30:@36827.4]
  assign _T_90913 = _T_90909[3]; // @[OneHot.scala 66:30:@36828.4]
  assign _T_90914 = _T_90909[4]; // @[OneHot.scala 66:30:@36829.4]
  assign _T_90915 = _T_90909[5]; // @[OneHot.scala 66:30:@36830.4]
  assign _T_90916 = _T_90909[6]; // @[OneHot.scala 66:30:@36831.4]
  assign _T_90917 = _T_90909[7]; // @[OneHot.scala 66:30:@36832.4]
  assign _T_90918 = _T_90909[8]; // @[OneHot.scala 66:30:@36833.4]
  assign _T_90919 = _T_90909[9]; // @[OneHot.scala 66:30:@36834.4]
  assign _T_90920 = _T_90909[10]; // @[OneHot.scala 66:30:@36835.4]
  assign _T_90921 = _T_90909[11]; // @[OneHot.scala 66:30:@36836.4]
  assign _T_90922 = _T_90909[12]; // @[OneHot.scala 66:30:@36837.4]
  assign _T_90923 = _T_90909[13]; // @[OneHot.scala 66:30:@36838.4]
  assign _T_90924 = _T_90909[14]; // @[OneHot.scala 66:30:@36839.4]
  assign _T_90925 = _T_90909[15]; // @[OneHot.scala 66:30:@36840.4]
  assign _T_90966 = loadRequest_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36858.4]
  assign _T_90967 = loadRequest_5 ? 16'h4000 : _T_90966; // @[Mux.scala 31:69:@36859.4]
  assign _T_90968 = loadRequest_4 ? 16'h2000 : _T_90967; // @[Mux.scala 31:69:@36860.4]
  assign _T_90969 = loadRequest_3 ? 16'h1000 : _T_90968; // @[Mux.scala 31:69:@36861.4]
  assign _T_90970 = loadRequest_2 ? 16'h800 : _T_90969; // @[Mux.scala 31:69:@36862.4]
  assign _T_90971 = loadRequest_1 ? 16'h400 : _T_90970; // @[Mux.scala 31:69:@36863.4]
  assign _T_90972 = loadRequest_0 ? 16'h200 : _T_90971; // @[Mux.scala 31:69:@36864.4]
  assign _T_90973 = loadRequest_15 ? 16'h100 : _T_90972; // @[Mux.scala 31:69:@36865.4]
  assign _T_90974 = loadRequest_14 ? 16'h80 : _T_90973; // @[Mux.scala 31:69:@36866.4]
  assign _T_90975 = loadRequest_13 ? 16'h40 : _T_90974; // @[Mux.scala 31:69:@36867.4]
  assign _T_90976 = loadRequest_12 ? 16'h20 : _T_90975; // @[Mux.scala 31:69:@36868.4]
  assign _T_90977 = loadRequest_11 ? 16'h10 : _T_90976; // @[Mux.scala 31:69:@36869.4]
  assign _T_90978 = loadRequest_10 ? 16'h8 : _T_90977; // @[Mux.scala 31:69:@36870.4]
  assign _T_90979 = loadRequest_9 ? 16'h4 : _T_90978; // @[Mux.scala 31:69:@36871.4]
  assign _T_90980 = loadRequest_8 ? 16'h2 : _T_90979; // @[Mux.scala 31:69:@36872.4]
  assign _T_90981 = loadRequest_7 ? 16'h1 : _T_90980; // @[Mux.scala 31:69:@36873.4]
  assign _T_90982 = _T_90981[0]; // @[OneHot.scala 66:30:@36874.4]
  assign _T_90983 = _T_90981[1]; // @[OneHot.scala 66:30:@36875.4]
  assign _T_90984 = _T_90981[2]; // @[OneHot.scala 66:30:@36876.4]
  assign _T_90985 = _T_90981[3]; // @[OneHot.scala 66:30:@36877.4]
  assign _T_90986 = _T_90981[4]; // @[OneHot.scala 66:30:@36878.4]
  assign _T_90987 = _T_90981[5]; // @[OneHot.scala 66:30:@36879.4]
  assign _T_90988 = _T_90981[6]; // @[OneHot.scala 66:30:@36880.4]
  assign _T_90989 = _T_90981[7]; // @[OneHot.scala 66:30:@36881.4]
  assign _T_90990 = _T_90981[8]; // @[OneHot.scala 66:30:@36882.4]
  assign _T_90991 = _T_90981[9]; // @[OneHot.scala 66:30:@36883.4]
  assign _T_90992 = _T_90981[10]; // @[OneHot.scala 66:30:@36884.4]
  assign _T_90993 = _T_90981[11]; // @[OneHot.scala 66:30:@36885.4]
  assign _T_90994 = _T_90981[12]; // @[OneHot.scala 66:30:@36886.4]
  assign _T_90995 = _T_90981[13]; // @[OneHot.scala 66:30:@36887.4]
  assign _T_90996 = _T_90981[14]; // @[OneHot.scala 66:30:@36888.4]
  assign _T_90997 = _T_90981[15]; // @[OneHot.scala 66:30:@36889.4]
  assign _T_91038 = loadRequest_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36907.4]
  assign _T_91039 = loadRequest_6 ? 16'h4000 : _T_91038; // @[Mux.scala 31:69:@36908.4]
  assign _T_91040 = loadRequest_5 ? 16'h2000 : _T_91039; // @[Mux.scala 31:69:@36909.4]
  assign _T_91041 = loadRequest_4 ? 16'h1000 : _T_91040; // @[Mux.scala 31:69:@36910.4]
  assign _T_91042 = loadRequest_3 ? 16'h800 : _T_91041; // @[Mux.scala 31:69:@36911.4]
  assign _T_91043 = loadRequest_2 ? 16'h400 : _T_91042; // @[Mux.scala 31:69:@36912.4]
  assign _T_91044 = loadRequest_1 ? 16'h200 : _T_91043; // @[Mux.scala 31:69:@36913.4]
  assign _T_91045 = loadRequest_0 ? 16'h100 : _T_91044; // @[Mux.scala 31:69:@36914.4]
  assign _T_91046 = loadRequest_15 ? 16'h80 : _T_91045; // @[Mux.scala 31:69:@36915.4]
  assign _T_91047 = loadRequest_14 ? 16'h40 : _T_91046; // @[Mux.scala 31:69:@36916.4]
  assign _T_91048 = loadRequest_13 ? 16'h20 : _T_91047; // @[Mux.scala 31:69:@36917.4]
  assign _T_91049 = loadRequest_12 ? 16'h10 : _T_91048; // @[Mux.scala 31:69:@36918.4]
  assign _T_91050 = loadRequest_11 ? 16'h8 : _T_91049; // @[Mux.scala 31:69:@36919.4]
  assign _T_91051 = loadRequest_10 ? 16'h4 : _T_91050; // @[Mux.scala 31:69:@36920.4]
  assign _T_91052 = loadRequest_9 ? 16'h2 : _T_91051; // @[Mux.scala 31:69:@36921.4]
  assign _T_91053 = loadRequest_8 ? 16'h1 : _T_91052; // @[Mux.scala 31:69:@36922.4]
  assign _T_91054 = _T_91053[0]; // @[OneHot.scala 66:30:@36923.4]
  assign _T_91055 = _T_91053[1]; // @[OneHot.scala 66:30:@36924.4]
  assign _T_91056 = _T_91053[2]; // @[OneHot.scala 66:30:@36925.4]
  assign _T_91057 = _T_91053[3]; // @[OneHot.scala 66:30:@36926.4]
  assign _T_91058 = _T_91053[4]; // @[OneHot.scala 66:30:@36927.4]
  assign _T_91059 = _T_91053[5]; // @[OneHot.scala 66:30:@36928.4]
  assign _T_91060 = _T_91053[6]; // @[OneHot.scala 66:30:@36929.4]
  assign _T_91061 = _T_91053[7]; // @[OneHot.scala 66:30:@36930.4]
  assign _T_91062 = _T_91053[8]; // @[OneHot.scala 66:30:@36931.4]
  assign _T_91063 = _T_91053[9]; // @[OneHot.scala 66:30:@36932.4]
  assign _T_91064 = _T_91053[10]; // @[OneHot.scala 66:30:@36933.4]
  assign _T_91065 = _T_91053[11]; // @[OneHot.scala 66:30:@36934.4]
  assign _T_91066 = _T_91053[12]; // @[OneHot.scala 66:30:@36935.4]
  assign _T_91067 = _T_91053[13]; // @[OneHot.scala 66:30:@36936.4]
  assign _T_91068 = _T_91053[14]; // @[OneHot.scala 66:30:@36937.4]
  assign _T_91069 = _T_91053[15]; // @[OneHot.scala 66:30:@36938.4]
  assign _T_91110 = loadRequest_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@36956.4]
  assign _T_91111 = loadRequest_7 ? 16'h4000 : _T_91110; // @[Mux.scala 31:69:@36957.4]
  assign _T_91112 = loadRequest_6 ? 16'h2000 : _T_91111; // @[Mux.scala 31:69:@36958.4]
  assign _T_91113 = loadRequest_5 ? 16'h1000 : _T_91112; // @[Mux.scala 31:69:@36959.4]
  assign _T_91114 = loadRequest_4 ? 16'h800 : _T_91113; // @[Mux.scala 31:69:@36960.4]
  assign _T_91115 = loadRequest_3 ? 16'h400 : _T_91114; // @[Mux.scala 31:69:@36961.4]
  assign _T_91116 = loadRequest_2 ? 16'h200 : _T_91115; // @[Mux.scala 31:69:@36962.4]
  assign _T_91117 = loadRequest_1 ? 16'h100 : _T_91116; // @[Mux.scala 31:69:@36963.4]
  assign _T_91118 = loadRequest_0 ? 16'h80 : _T_91117; // @[Mux.scala 31:69:@36964.4]
  assign _T_91119 = loadRequest_15 ? 16'h40 : _T_91118; // @[Mux.scala 31:69:@36965.4]
  assign _T_91120 = loadRequest_14 ? 16'h20 : _T_91119; // @[Mux.scala 31:69:@36966.4]
  assign _T_91121 = loadRequest_13 ? 16'h10 : _T_91120; // @[Mux.scala 31:69:@36967.4]
  assign _T_91122 = loadRequest_12 ? 16'h8 : _T_91121; // @[Mux.scala 31:69:@36968.4]
  assign _T_91123 = loadRequest_11 ? 16'h4 : _T_91122; // @[Mux.scala 31:69:@36969.4]
  assign _T_91124 = loadRequest_10 ? 16'h2 : _T_91123; // @[Mux.scala 31:69:@36970.4]
  assign _T_91125 = loadRequest_9 ? 16'h1 : _T_91124; // @[Mux.scala 31:69:@36971.4]
  assign _T_91126 = _T_91125[0]; // @[OneHot.scala 66:30:@36972.4]
  assign _T_91127 = _T_91125[1]; // @[OneHot.scala 66:30:@36973.4]
  assign _T_91128 = _T_91125[2]; // @[OneHot.scala 66:30:@36974.4]
  assign _T_91129 = _T_91125[3]; // @[OneHot.scala 66:30:@36975.4]
  assign _T_91130 = _T_91125[4]; // @[OneHot.scala 66:30:@36976.4]
  assign _T_91131 = _T_91125[5]; // @[OneHot.scala 66:30:@36977.4]
  assign _T_91132 = _T_91125[6]; // @[OneHot.scala 66:30:@36978.4]
  assign _T_91133 = _T_91125[7]; // @[OneHot.scala 66:30:@36979.4]
  assign _T_91134 = _T_91125[8]; // @[OneHot.scala 66:30:@36980.4]
  assign _T_91135 = _T_91125[9]; // @[OneHot.scala 66:30:@36981.4]
  assign _T_91136 = _T_91125[10]; // @[OneHot.scala 66:30:@36982.4]
  assign _T_91137 = _T_91125[11]; // @[OneHot.scala 66:30:@36983.4]
  assign _T_91138 = _T_91125[12]; // @[OneHot.scala 66:30:@36984.4]
  assign _T_91139 = _T_91125[13]; // @[OneHot.scala 66:30:@36985.4]
  assign _T_91140 = _T_91125[14]; // @[OneHot.scala 66:30:@36986.4]
  assign _T_91141 = _T_91125[15]; // @[OneHot.scala 66:30:@36987.4]
  assign _T_91182 = loadRequest_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37005.4]
  assign _T_91183 = loadRequest_8 ? 16'h4000 : _T_91182; // @[Mux.scala 31:69:@37006.4]
  assign _T_91184 = loadRequest_7 ? 16'h2000 : _T_91183; // @[Mux.scala 31:69:@37007.4]
  assign _T_91185 = loadRequest_6 ? 16'h1000 : _T_91184; // @[Mux.scala 31:69:@37008.4]
  assign _T_91186 = loadRequest_5 ? 16'h800 : _T_91185; // @[Mux.scala 31:69:@37009.4]
  assign _T_91187 = loadRequest_4 ? 16'h400 : _T_91186; // @[Mux.scala 31:69:@37010.4]
  assign _T_91188 = loadRequest_3 ? 16'h200 : _T_91187; // @[Mux.scala 31:69:@37011.4]
  assign _T_91189 = loadRequest_2 ? 16'h100 : _T_91188; // @[Mux.scala 31:69:@37012.4]
  assign _T_91190 = loadRequest_1 ? 16'h80 : _T_91189; // @[Mux.scala 31:69:@37013.4]
  assign _T_91191 = loadRequest_0 ? 16'h40 : _T_91190; // @[Mux.scala 31:69:@37014.4]
  assign _T_91192 = loadRequest_15 ? 16'h20 : _T_91191; // @[Mux.scala 31:69:@37015.4]
  assign _T_91193 = loadRequest_14 ? 16'h10 : _T_91192; // @[Mux.scala 31:69:@37016.4]
  assign _T_91194 = loadRequest_13 ? 16'h8 : _T_91193; // @[Mux.scala 31:69:@37017.4]
  assign _T_91195 = loadRequest_12 ? 16'h4 : _T_91194; // @[Mux.scala 31:69:@37018.4]
  assign _T_91196 = loadRequest_11 ? 16'h2 : _T_91195; // @[Mux.scala 31:69:@37019.4]
  assign _T_91197 = loadRequest_10 ? 16'h1 : _T_91196; // @[Mux.scala 31:69:@37020.4]
  assign _T_91198 = _T_91197[0]; // @[OneHot.scala 66:30:@37021.4]
  assign _T_91199 = _T_91197[1]; // @[OneHot.scala 66:30:@37022.4]
  assign _T_91200 = _T_91197[2]; // @[OneHot.scala 66:30:@37023.4]
  assign _T_91201 = _T_91197[3]; // @[OneHot.scala 66:30:@37024.4]
  assign _T_91202 = _T_91197[4]; // @[OneHot.scala 66:30:@37025.4]
  assign _T_91203 = _T_91197[5]; // @[OneHot.scala 66:30:@37026.4]
  assign _T_91204 = _T_91197[6]; // @[OneHot.scala 66:30:@37027.4]
  assign _T_91205 = _T_91197[7]; // @[OneHot.scala 66:30:@37028.4]
  assign _T_91206 = _T_91197[8]; // @[OneHot.scala 66:30:@37029.4]
  assign _T_91207 = _T_91197[9]; // @[OneHot.scala 66:30:@37030.4]
  assign _T_91208 = _T_91197[10]; // @[OneHot.scala 66:30:@37031.4]
  assign _T_91209 = _T_91197[11]; // @[OneHot.scala 66:30:@37032.4]
  assign _T_91210 = _T_91197[12]; // @[OneHot.scala 66:30:@37033.4]
  assign _T_91211 = _T_91197[13]; // @[OneHot.scala 66:30:@37034.4]
  assign _T_91212 = _T_91197[14]; // @[OneHot.scala 66:30:@37035.4]
  assign _T_91213 = _T_91197[15]; // @[OneHot.scala 66:30:@37036.4]
  assign _T_91254 = loadRequest_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37054.4]
  assign _T_91255 = loadRequest_9 ? 16'h4000 : _T_91254; // @[Mux.scala 31:69:@37055.4]
  assign _T_91256 = loadRequest_8 ? 16'h2000 : _T_91255; // @[Mux.scala 31:69:@37056.4]
  assign _T_91257 = loadRequest_7 ? 16'h1000 : _T_91256; // @[Mux.scala 31:69:@37057.4]
  assign _T_91258 = loadRequest_6 ? 16'h800 : _T_91257; // @[Mux.scala 31:69:@37058.4]
  assign _T_91259 = loadRequest_5 ? 16'h400 : _T_91258; // @[Mux.scala 31:69:@37059.4]
  assign _T_91260 = loadRequest_4 ? 16'h200 : _T_91259; // @[Mux.scala 31:69:@37060.4]
  assign _T_91261 = loadRequest_3 ? 16'h100 : _T_91260; // @[Mux.scala 31:69:@37061.4]
  assign _T_91262 = loadRequest_2 ? 16'h80 : _T_91261; // @[Mux.scala 31:69:@37062.4]
  assign _T_91263 = loadRequest_1 ? 16'h40 : _T_91262; // @[Mux.scala 31:69:@37063.4]
  assign _T_91264 = loadRequest_0 ? 16'h20 : _T_91263; // @[Mux.scala 31:69:@37064.4]
  assign _T_91265 = loadRequest_15 ? 16'h10 : _T_91264; // @[Mux.scala 31:69:@37065.4]
  assign _T_91266 = loadRequest_14 ? 16'h8 : _T_91265; // @[Mux.scala 31:69:@37066.4]
  assign _T_91267 = loadRequest_13 ? 16'h4 : _T_91266; // @[Mux.scala 31:69:@37067.4]
  assign _T_91268 = loadRequest_12 ? 16'h2 : _T_91267; // @[Mux.scala 31:69:@37068.4]
  assign _T_91269 = loadRequest_11 ? 16'h1 : _T_91268; // @[Mux.scala 31:69:@37069.4]
  assign _T_91270 = _T_91269[0]; // @[OneHot.scala 66:30:@37070.4]
  assign _T_91271 = _T_91269[1]; // @[OneHot.scala 66:30:@37071.4]
  assign _T_91272 = _T_91269[2]; // @[OneHot.scala 66:30:@37072.4]
  assign _T_91273 = _T_91269[3]; // @[OneHot.scala 66:30:@37073.4]
  assign _T_91274 = _T_91269[4]; // @[OneHot.scala 66:30:@37074.4]
  assign _T_91275 = _T_91269[5]; // @[OneHot.scala 66:30:@37075.4]
  assign _T_91276 = _T_91269[6]; // @[OneHot.scala 66:30:@37076.4]
  assign _T_91277 = _T_91269[7]; // @[OneHot.scala 66:30:@37077.4]
  assign _T_91278 = _T_91269[8]; // @[OneHot.scala 66:30:@37078.4]
  assign _T_91279 = _T_91269[9]; // @[OneHot.scala 66:30:@37079.4]
  assign _T_91280 = _T_91269[10]; // @[OneHot.scala 66:30:@37080.4]
  assign _T_91281 = _T_91269[11]; // @[OneHot.scala 66:30:@37081.4]
  assign _T_91282 = _T_91269[12]; // @[OneHot.scala 66:30:@37082.4]
  assign _T_91283 = _T_91269[13]; // @[OneHot.scala 66:30:@37083.4]
  assign _T_91284 = _T_91269[14]; // @[OneHot.scala 66:30:@37084.4]
  assign _T_91285 = _T_91269[15]; // @[OneHot.scala 66:30:@37085.4]
  assign _T_91326 = loadRequest_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37103.4]
  assign _T_91327 = loadRequest_10 ? 16'h4000 : _T_91326; // @[Mux.scala 31:69:@37104.4]
  assign _T_91328 = loadRequest_9 ? 16'h2000 : _T_91327; // @[Mux.scala 31:69:@37105.4]
  assign _T_91329 = loadRequest_8 ? 16'h1000 : _T_91328; // @[Mux.scala 31:69:@37106.4]
  assign _T_91330 = loadRequest_7 ? 16'h800 : _T_91329; // @[Mux.scala 31:69:@37107.4]
  assign _T_91331 = loadRequest_6 ? 16'h400 : _T_91330; // @[Mux.scala 31:69:@37108.4]
  assign _T_91332 = loadRequest_5 ? 16'h200 : _T_91331; // @[Mux.scala 31:69:@37109.4]
  assign _T_91333 = loadRequest_4 ? 16'h100 : _T_91332; // @[Mux.scala 31:69:@37110.4]
  assign _T_91334 = loadRequest_3 ? 16'h80 : _T_91333; // @[Mux.scala 31:69:@37111.4]
  assign _T_91335 = loadRequest_2 ? 16'h40 : _T_91334; // @[Mux.scala 31:69:@37112.4]
  assign _T_91336 = loadRequest_1 ? 16'h20 : _T_91335; // @[Mux.scala 31:69:@37113.4]
  assign _T_91337 = loadRequest_0 ? 16'h10 : _T_91336; // @[Mux.scala 31:69:@37114.4]
  assign _T_91338 = loadRequest_15 ? 16'h8 : _T_91337; // @[Mux.scala 31:69:@37115.4]
  assign _T_91339 = loadRequest_14 ? 16'h4 : _T_91338; // @[Mux.scala 31:69:@37116.4]
  assign _T_91340 = loadRequest_13 ? 16'h2 : _T_91339; // @[Mux.scala 31:69:@37117.4]
  assign _T_91341 = loadRequest_12 ? 16'h1 : _T_91340; // @[Mux.scala 31:69:@37118.4]
  assign _T_91342 = _T_91341[0]; // @[OneHot.scala 66:30:@37119.4]
  assign _T_91343 = _T_91341[1]; // @[OneHot.scala 66:30:@37120.4]
  assign _T_91344 = _T_91341[2]; // @[OneHot.scala 66:30:@37121.4]
  assign _T_91345 = _T_91341[3]; // @[OneHot.scala 66:30:@37122.4]
  assign _T_91346 = _T_91341[4]; // @[OneHot.scala 66:30:@37123.4]
  assign _T_91347 = _T_91341[5]; // @[OneHot.scala 66:30:@37124.4]
  assign _T_91348 = _T_91341[6]; // @[OneHot.scala 66:30:@37125.4]
  assign _T_91349 = _T_91341[7]; // @[OneHot.scala 66:30:@37126.4]
  assign _T_91350 = _T_91341[8]; // @[OneHot.scala 66:30:@37127.4]
  assign _T_91351 = _T_91341[9]; // @[OneHot.scala 66:30:@37128.4]
  assign _T_91352 = _T_91341[10]; // @[OneHot.scala 66:30:@37129.4]
  assign _T_91353 = _T_91341[11]; // @[OneHot.scala 66:30:@37130.4]
  assign _T_91354 = _T_91341[12]; // @[OneHot.scala 66:30:@37131.4]
  assign _T_91355 = _T_91341[13]; // @[OneHot.scala 66:30:@37132.4]
  assign _T_91356 = _T_91341[14]; // @[OneHot.scala 66:30:@37133.4]
  assign _T_91357 = _T_91341[15]; // @[OneHot.scala 66:30:@37134.4]
  assign _T_91398 = loadRequest_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37152.4]
  assign _T_91399 = loadRequest_11 ? 16'h4000 : _T_91398; // @[Mux.scala 31:69:@37153.4]
  assign _T_91400 = loadRequest_10 ? 16'h2000 : _T_91399; // @[Mux.scala 31:69:@37154.4]
  assign _T_91401 = loadRequest_9 ? 16'h1000 : _T_91400; // @[Mux.scala 31:69:@37155.4]
  assign _T_91402 = loadRequest_8 ? 16'h800 : _T_91401; // @[Mux.scala 31:69:@37156.4]
  assign _T_91403 = loadRequest_7 ? 16'h400 : _T_91402; // @[Mux.scala 31:69:@37157.4]
  assign _T_91404 = loadRequest_6 ? 16'h200 : _T_91403; // @[Mux.scala 31:69:@37158.4]
  assign _T_91405 = loadRequest_5 ? 16'h100 : _T_91404; // @[Mux.scala 31:69:@37159.4]
  assign _T_91406 = loadRequest_4 ? 16'h80 : _T_91405; // @[Mux.scala 31:69:@37160.4]
  assign _T_91407 = loadRequest_3 ? 16'h40 : _T_91406; // @[Mux.scala 31:69:@37161.4]
  assign _T_91408 = loadRequest_2 ? 16'h20 : _T_91407; // @[Mux.scala 31:69:@37162.4]
  assign _T_91409 = loadRequest_1 ? 16'h10 : _T_91408; // @[Mux.scala 31:69:@37163.4]
  assign _T_91410 = loadRequest_0 ? 16'h8 : _T_91409; // @[Mux.scala 31:69:@37164.4]
  assign _T_91411 = loadRequest_15 ? 16'h4 : _T_91410; // @[Mux.scala 31:69:@37165.4]
  assign _T_91412 = loadRequest_14 ? 16'h2 : _T_91411; // @[Mux.scala 31:69:@37166.4]
  assign _T_91413 = loadRequest_13 ? 16'h1 : _T_91412; // @[Mux.scala 31:69:@37167.4]
  assign _T_91414 = _T_91413[0]; // @[OneHot.scala 66:30:@37168.4]
  assign _T_91415 = _T_91413[1]; // @[OneHot.scala 66:30:@37169.4]
  assign _T_91416 = _T_91413[2]; // @[OneHot.scala 66:30:@37170.4]
  assign _T_91417 = _T_91413[3]; // @[OneHot.scala 66:30:@37171.4]
  assign _T_91418 = _T_91413[4]; // @[OneHot.scala 66:30:@37172.4]
  assign _T_91419 = _T_91413[5]; // @[OneHot.scala 66:30:@37173.4]
  assign _T_91420 = _T_91413[6]; // @[OneHot.scala 66:30:@37174.4]
  assign _T_91421 = _T_91413[7]; // @[OneHot.scala 66:30:@37175.4]
  assign _T_91422 = _T_91413[8]; // @[OneHot.scala 66:30:@37176.4]
  assign _T_91423 = _T_91413[9]; // @[OneHot.scala 66:30:@37177.4]
  assign _T_91424 = _T_91413[10]; // @[OneHot.scala 66:30:@37178.4]
  assign _T_91425 = _T_91413[11]; // @[OneHot.scala 66:30:@37179.4]
  assign _T_91426 = _T_91413[12]; // @[OneHot.scala 66:30:@37180.4]
  assign _T_91427 = _T_91413[13]; // @[OneHot.scala 66:30:@37181.4]
  assign _T_91428 = _T_91413[14]; // @[OneHot.scala 66:30:@37182.4]
  assign _T_91429 = _T_91413[15]; // @[OneHot.scala 66:30:@37183.4]
  assign _T_91470 = loadRequest_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37201.4]
  assign _T_91471 = loadRequest_12 ? 16'h4000 : _T_91470; // @[Mux.scala 31:69:@37202.4]
  assign _T_91472 = loadRequest_11 ? 16'h2000 : _T_91471; // @[Mux.scala 31:69:@37203.4]
  assign _T_91473 = loadRequest_10 ? 16'h1000 : _T_91472; // @[Mux.scala 31:69:@37204.4]
  assign _T_91474 = loadRequest_9 ? 16'h800 : _T_91473; // @[Mux.scala 31:69:@37205.4]
  assign _T_91475 = loadRequest_8 ? 16'h400 : _T_91474; // @[Mux.scala 31:69:@37206.4]
  assign _T_91476 = loadRequest_7 ? 16'h200 : _T_91475; // @[Mux.scala 31:69:@37207.4]
  assign _T_91477 = loadRequest_6 ? 16'h100 : _T_91476; // @[Mux.scala 31:69:@37208.4]
  assign _T_91478 = loadRequest_5 ? 16'h80 : _T_91477; // @[Mux.scala 31:69:@37209.4]
  assign _T_91479 = loadRequest_4 ? 16'h40 : _T_91478; // @[Mux.scala 31:69:@37210.4]
  assign _T_91480 = loadRequest_3 ? 16'h20 : _T_91479; // @[Mux.scala 31:69:@37211.4]
  assign _T_91481 = loadRequest_2 ? 16'h10 : _T_91480; // @[Mux.scala 31:69:@37212.4]
  assign _T_91482 = loadRequest_1 ? 16'h8 : _T_91481; // @[Mux.scala 31:69:@37213.4]
  assign _T_91483 = loadRequest_0 ? 16'h4 : _T_91482; // @[Mux.scala 31:69:@37214.4]
  assign _T_91484 = loadRequest_15 ? 16'h2 : _T_91483; // @[Mux.scala 31:69:@37215.4]
  assign _T_91485 = loadRequest_14 ? 16'h1 : _T_91484; // @[Mux.scala 31:69:@37216.4]
  assign _T_91486 = _T_91485[0]; // @[OneHot.scala 66:30:@37217.4]
  assign _T_91487 = _T_91485[1]; // @[OneHot.scala 66:30:@37218.4]
  assign _T_91488 = _T_91485[2]; // @[OneHot.scala 66:30:@37219.4]
  assign _T_91489 = _T_91485[3]; // @[OneHot.scala 66:30:@37220.4]
  assign _T_91490 = _T_91485[4]; // @[OneHot.scala 66:30:@37221.4]
  assign _T_91491 = _T_91485[5]; // @[OneHot.scala 66:30:@37222.4]
  assign _T_91492 = _T_91485[6]; // @[OneHot.scala 66:30:@37223.4]
  assign _T_91493 = _T_91485[7]; // @[OneHot.scala 66:30:@37224.4]
  assign _T_91494 = _T_91485[8]; // @[OneHot.scala 66:30:@37225.4]
  assign _T_91495 = _T_91485[9]; // @[OneHot.scala 66:30:@37226.4]
  assign _T_91496 = _T_91485[10]; // @[OneHot.scala 66:30:@37227.4]
  assign _T_91497 = _T_91485[11]; // @[OneHot.scala 66:30:@37228.4]
  assign _T_91498 = _T_91485[12]; // @[OneHot.scala 66:30:@37229.4]
  assign _T_91499 = _T_91485[13]; // @[OneHot.scala 66:30:@37230.4]
  assign _T_91500 = _T_91485[14]; // @[OneHot.scala 66:30:@37231.4]
  assign _T_91501 = _T_91485[15]; // @[OneHot.scala 66:30:@37232.4]
  assign _T_91542 = loadRequest_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@37250.4]
  assign _T_91543 = loadRequest_13 ? 16'h4000 : _T_91542; // @[Mux.scala 31:69:@37251.4]
  assign _T_91544 = loadRequest_12 ? 16'h2000 : _T_91543; // @[Mux.scala 31:69:@37252.4]
  assign _T_91545 = loadRequest_11 ? 16'h1000 : _T_91544; // @[Mux.scala 31:69:@37253.4]
  assign _T_91546 = loadRequest_10 ? 16'h800 : _T_91545; // @[Mux.scala 31:69:@37254.4]
  assign _T_91547 = loadRequest_9 ? 16'h400 : _T_91546; // @[Mux.scala 31:69:@37255.4]
  assign _T_91548 = loadRequest_8 ? 16'h200 : _T_91547; // @[Mux.scala 31:69:@37256.4]
  assign _T_91549 = loadRequest_7 ? 16'h100 : _T_91548; // @[Mux.scala 31:69:@37257.4]
  assign _T_91550 = loadRequest_6 ? 16'h80 : _T_91549; // @[Mux.scala 31:69:@37258.4]
  assign _T_91551 = loadRequest_5 ? 16'h40 : _T_91550; // @[Mux.scala 31:69:@37259.4]
  assign _T_91552 = loadRequest_4 ? 16'h20 : _T_91551; // @[Mux.scala 31:69:@37260.4]
  assign _T_91553 = loadRequest_3 ? 16'h10 : _T_91552; // @[Mux.scala 31:69:@37261.4]
  assign _T_91554 = loadRequest_2 ? 16'h8 : _T_91553; // @[Mux.scala 31:69:@37262.4]
  assign _T_91555 = loadRequest_1 ? 16'h4 : _T_91554; // @[Mux.scala 31:69:@37263.4]
  assign _T_91556 = loadRequest_0 ? 16'h2 : _T_91555; // @[Mux.scala 31:69:@37264.4]
  assign _T_91557 = loadRequest_15 ? 16'h1 : _T_91556; // @[Mux.scala 31:69:@37265.4]
  assign _T_91558 = _T_91557[0]; // @[OneHot.scala 66:30:@37266.4]
  assign _T_91559 = _T_91557[1]; // @[OneHot.scala 66:30:@37267.4]
  assign _T_91560 = _T_91557[2]; // @[OneHot.scala 66:30:@37268.4]
  assign _T_91561 = _T_91557[3]; // @[OneHot.scala 66:30:@37269.4]
  assign _T_91562 = _T_91557[4]; // @[OneHot.scala 66:30:@37270.4]
  assign _T_91563 = _T_91557[5]; // @[OneHot.scala 66:30:@37271.4]
  assign _T_91564 = _T_91557[6]; // @[OneHot.scala 66:30:@37272.4]
  assign _T_91565 = _T_91557[7]; // @[OneHot.scala 66:30:@37273.4]
  assign _T_91566 = _T_91557[8]; // @[OneHot.scala 66:30:@37274.4]
  assign _T_91567 = _T_91557[9]; // @[OneHot.scala 66:30:@37275.4]
  assign _T_91568 = _T_91557[10]; // @[OneHot.scala 66:30:@37276.4]
  assign _T_91569 = _T_91557[11]; // @[OneHot.scala 66:30:@37277.4]
  assign _T_91570 = _T_91557[12]; // @[OneHot.scala 66:30:@37278.4]
  assign _T_91571 = _T_91557[13]; // @[OneHot.scala 66:30:@37279.4]
  assign _T_91572 = _T_91557[14]; // @[OneHot.scala 66:30:@37280.4]
  assign _T_91573 = _T_91557[15]; // @[OneHot.scala 66:30:@37281.4]
  assign _T_91638 = {_T_90485,_T_90484,_T_90483,_T_90482,_T_90481,_T_90480,_T_90479,_T_90478}; // @[Mux.scala 19:72:@37305.4]
  assign _T_91646 = {_T_90493,_T_90492,_T_90491,_T_90490,_T_90489,_T_90488,_T_90487,_T_90486,_T_91638}; // @[Mux.scala 19:72:@37313.4]
  assign _T_91648 = _T_90406 ? _T_91646 : 16'h0; // @[Mux.scala 19:72:@37314.4]
  assign _T_91655 = {_T_90556,_T_90555,_T_90554,_T_90553,_T_90552,_T_90551,_T_90550,_T_90565}; // @[Mux.scala 19:72:@37321.4]
  assign _T_91663 = {_T_90564,_T_90563,_T_90562,_T_90561,_T_90560,_T_90559,_T_90558,_T_90557,_T_91655}; // @[Mux.scala 19:72:@37329.4]
  assign _T_91665 = _T_90407 ? _T_91663 : 16'h0; // @[Mux.scala 19:72:@37330.4]
  assign _T_91672 = {_T_90627,_T_90626,_T_90625,_T_90624,_T_90623,_T_90622,_T_90637,_T_90636}; // @[Mux.scala 19:72:@37337.4]
  assign _T_91680 = {_T_90635,_T_90634,_T_90633,_T_90632,_T_90631,_T_90630,_T_90629,_T_90628,_T_91672}; // @[Mux.scala 19:72:@37345.4]
  assign _T_91682 = _T_90408 ? _T_91680 : 16'h0; // @[Mux.scala 19:72:@37346.4]
  assign _T_91689 = {_T_90698,_T_90697,_T_90696,_T_90695,_T_90694,_T_90709,_T_90708,_T_90707}; // @[Mux.scala 19:72:@37353.4]
  assign _T_91697 = {_T_90706,_T_90705,_T_90704,_T_90703,_T_90702,_T_90701,_T_90700,_T_90699,_T_91689}; // @[Mux.scala 19:72:@37361.4]
  assign _T_91699 = _T_90409 ? _T_91697 : 16'h0; // @[Mux.scala 19:72:@37362.4]
  assign _T_91706 = {_T_90769,_T_90768,_T_90767,_T_90766,_T_90781,_T_90780,_T_90779,_T_90778}; // @[Mux.scala 19:72:@37369.4]
  assign _T_91714 = {_T_90777,_T_90776,_T_90775,_T_90774,_T_90773,_T_90772,_T_90771,_T_90770,_T_91706}; // @[Mux.scala 19:72:@37377.4]
  assign _T_91716 = _T_90410 ? _T_91714 : 16'h0; // @[Mux.scala 19:72:@37378.4]
  assign _T_91723 = {_T_90840,_T_90839,_T_90838,_T_90853,_T_90852,_T_90851,_T_90850,_T_90849}; // @[Mux.scala 19:72:@37385.4]
  assign _T_91731 = {_T_90848,_T_90847,_T_90846,_T_90845,_T_90844,_T_90843,_T_90842,_T_90841,_T_91723}; // @[Mux.scala 19:72:@37393.4]
  assign _T_91733 = _T_90411 ? _T_91731 : 16'h0; // @[Mux.scala 19:72:@37394.4]
  assign _T_91740 = {_T_90911,_T_90910,_T_90925,_T_90924,_T_90923,_T_90922,_T_90921,_T_90920}; // @[Mux.scala 19:72:@37401.4]
  assign _T_91748 = {_T_90919,_T_90918,_T_90917,_T_90916,_T_90915,_T_90914,_T_90913,_T_90912,_T_91740}; // @[Mux.scala 19:72:@37409.4]
  assign _T_91750 = _T_90412 ? _T_91748 : 16'h0; // @[Mux.scala 19:72:@37410.4]
  assign _T_91757 = {_T_90982,_T_90997,_T_90996,_T_90995,_T_90994,_T_90993,_T_90992,_T_90991}; // @[Mux.scala 19:72:@37417.4]
  assign _T_91765 = {_T_90990,_T_90989,_T_90988,_T_90987,_T_90986,_T_90985,_T_90984,_T_90983,_T_91757}; // @[Mux.scala 19:72:@37425.4]
  assign _T_91767 = _T_90413 ? _T_91765 : 16'h0; // @[Mux.scala 19:72:@37426.4]
  assign _T_91774 = {_T_91069,_T_91068,_T_91067,_T_91066,_T_91065,_T_91064,_T_91063,_T_91062}; // @[Mux.scala 19:72:@37433.4]
  assign _T_91782 = {_T_91061,_T_91060,_T_91059,_T_91058,_T_91057,_T_91056,_T_91055,_T_91054,_T_91774}; // @[Mux.scala 19:72:@37441.4]
  assign _T_91784 = _T_90414 ? _T_91782 : 16'h0; // @[Mux.scala 19:72:@37442.4]
  assign _T_91791 = {_T_91140,_T_91139,_T_91138,_T_91137,_T_91136,_T_91135,_T_91134,_T_91133}; // @[Mux.scala 19:72:@37449.4]
  assign _T_91799 = {_T_91132,_T_91131,_T_91130,_T_91129,_T_91128,_T_91127,_T_91126,_T_91141,_T_91791}; // @[Mux.scala 19:72:@37457.4]
  assign _T_91801 = _T_90415 ? _T_91799 : 16'h0; // @[Mux.scala 19:72:@37458.4]
  assign _T_91808 = {_T_91211,_T_91210,_T_91209,_T_91208,_T_91207,_T_91206,_T_91205,_T_91204}; // @[Mux.scala 19:72:@37465.4]
  assign _T_91816 = {_T_91203,_T_91202,_T_91201,_T_91200,_T_91199,_T_91198,_T_91213,_T_91212,_T_91808}; // @[Mux.scala 19:72:@37473.4]
  assign _T_91818 = _T_90416 ? _T_91816 : 16'h0; // @[Mux.scala 19:72:@37474.4]
  assign _T_91825 = {_T_91282,_T_91281,_T_91280,_T_91279,_T_91278,_T_91277,_T_91276,_T_91275}; // @[Mux.scala 19:72:@37481.4]
  assign _T_91833 = {_T_91274,_T_91273,_T_91272,_T_91271,_T_91270,_T_91285,_T_91284,_T_91283,_T_91825}; // @[Mux.scala 19:72:@37489.4]
  assign _T_91835 = _T_90417 ? _T_91833 : 16'h0; // @[Mux.scala 19:72:@37490.4]
  assign _T_91842 = {_T_91353,_T_91352,_T_91351,_T_91350,_T_91349,_T_91348,_T_91347,_T_91346}; // @[Mux.scala 19:72:@37497.4]
  assign _T_91850 = {_T_91345,_T_91344,_T_91343,_T_91342,_T_91357,_T_91356,_T_91355,_T_91354,_T_91842}; // @[Mux.scala 19:72:@37505.4]
  assign _T_91852 = _T_90418 ? _T_91850 : 16'h0; // @[Mux.scala 19:72:@37506.4]
  assign _T_91859 = {_T_91424,_T_91423,_T_91422,_T_91421,_T_91420,_T_91419,_T_91418,_T_91417}; // @[Mux.scala 19:72:@37513.4]
  assign _T_91867 = {_T_91416,_T_91415,_T_91414,_T_91429,_T_91428,_T_91427,_T_91426,_T_91425,_T_91859}; // @[Mux.scala 19:72:@37521.4]
  assign _T_91869 = _T_90419 ? _T_91867 : 16'h0; // @[Mux.scala 19:72:@37522.4]
  assign _T_91876 = {_T_91495,_T_91494,_T_91493,_T_91492,_T_91491,_T_91490,_T_91489,_T_91488}; // @[Mux.scala 19:72:@37529.4]
  assign _T_91884 = {_T_91487,_T_91486,_T_91501,_T_91500,_T_91499,_T_91498,_T_91497,_T_91496,_T_91876}; // @[Mux.scala 19:72:@37537.4]
  assign _T_91886 = _T_90420 ? _T_91884 : 16'h0; // @[Mux.scala 19:72:@37538.4]
  assign _T_91893 = {_T_91566,_T_91565,_T_91564,_T_91563,_T_91562,_T_91561,_T_91560,_T_91559}; // @[Mux.scala 19:72:@37545.4]
  assign _T_91901 = {_T_91558,_T_91573,_T_91572,_T_91571,_T_91570,_T_91569,_T_91568,_T_91567,_T_91893}; // @[Mux.scala 19:72:@37553.4]
  assign _T_91903 = _T_90421 ? _T_91901 : 16'h0; // @[Mux.scala 19:72:@37554.4]
  assign _T_91904 = _T_91648 | _T_91665; // @[Mux.scala 19:72:@37555.4]
  assign _T_91905 = _T_91904 | _T_91682; // @[Mux.scala 19:72:@37556.4]
  assign _T_91906 = _T_91905 | _T_91699; // @[Mux.scala 19:72:@37557.4]
  assign _T_91907 = _T_91906 | _T_91716; // @[Mux.scala 19:72:@37558.4]
  assign _T_91908 = _T_91907 | _T_91733; // @[Mux.scala 19:72:@37559.4]
  assign _T_91909 = _T_91908 | _T_91750; // @[Mux.scala 19:72:@37560.4]
  assign _T_91910 = _T_91909 | _T_91767; // @[Mux.scala 19:72:@37561.4]
  assign _T_91911 = _T_91910 | _T_91784; // @[Mux.scala 19:72:@37562.4]
  assign _T_91912 = _T_91911 | _T_91801; // @[Mux.scala 19:72:@37563.4]
  assign _T_91913 = _T_91912 | _T_91818; // @[Mux.scala 19:72:@37564.4]
  assign _T_91914 = _T_91913 | _T_91835; // @[Mux.scala 19:72:@37565.4]
  assign _T_91915 = _T_91914 | _T_91852; // @[Mux.scala 19:72:@37566.4]
  assign _T_91916 = _T_91915 | _T_91869; // @[Mux.scala 19:72:@37567.4]
  assign _T_91917 = _T_91916 | _T_91886; // @[Mux.scala 19:72:@37568.4]
  assign _T_91918 = _T_91917 | _T_91903; // @[Mux.scala 19:72:@37569.4]
  assign priorityLoadRequest_0 = _T_91918[0]; // @[Mux.scala 19:72:@37573.4]
  assign priorityLoadRequest_1 = _T_91918[1]; // @[Mux.scala 19:72:@37575.4]
  assign priorityLoadRequest_2 = _T_91918[2]; // @[Mux.scala 19:72:@37577.4]
  assign priorityLoadRequest_3 = _T_91918[3]; // @[Mux.scala 19:72:@37579.4]
  assign priorityLoadRequest_4 = _T_91918[4]; // @[Mux.scala 19:72:@37581.4]
  assign priorityLoadRequest_5 = _T_91918[5]; // @[Mux.scala 19:72:@37583.4]
  assign priorityLoadRequest_6 = _T_91918[6]; // @[Mux.scala 19:72:@37585.4]
  assign priorityLoadRequest_7 = _T_91918[7]; // @[Mux.scala 19:72:@37587.4]
  assign priorityLoadRequest_8 = _T_91918[8]; // @[Mux.scala 19:72:@37589.4]
  assign priorityLoadRequest_9 = _T_91918[9]; // @[Mux.scala 19:72:@37591.4]
  assign priorityLoadRequest_10 = _T_91918[10]; // @[Mux.scala 19:72:@37593.4]
  assign priorityLoadRequest_11 = _T_91918[11]; // @[Mux.scala 19:72:@37595.4]
  assign priorityLoadRequest_12 = _T_91918[12]; // @[Mux.scala 19:72:@37597.4]
  assign priorityLoadRequest_13 = _T_91918[13]; // @[Mux.scala 19:72:@37599.4]
  assign priorityLoadRequest_14 = _T_91918[14]; // @[Mux.scala 19:72:@37601.4]
  assign priorityLoadRequest_15 = _T_91918[15]; // @[Mux.scala 19:72:@37603.4]
  assign _T_92186 = priorityLoadRequest_0 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37627.6]
  assign _GEN_1920 = _T_92186 ? 1'h1 : loadInitiated_0; // @[AxiLoadQueue.scala 212:70:@37628.6]
  assign _GEN_1921 = initBits_0 ? 1'h0 : _GEN_1920; // @[AxiLoadQueue.scala 210:22:@37623.4]
  assign _T_92189 = priorityLoadRequest_1 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37635.6]
  assign _GEN_1922 = _T_92189 ? 1'h1 : loadInitiated_1; // @[AxiLoadQueue.scala 212:70:@37636.6]
  assign _GEN_1923 = initBits_1 ? 1'h0 : _GEN_1922; // @[AxiLoadQueue.scala 210:22:@37631.4]
  assign _T_92192 = priorityLoadRequest_2 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37643.6]
  assign _GEN_1924 = _T_92192 ? 1'h1 : loadInitiated_2; // @[AxiLoadQueue.scala 212:70:@37644.6]
  assign _GEN_1925 = initBits_2 ? 1'h0 : _GEN_1924; // @[AxiLoadQueue.scala 210:22:@37639.4]
  assign _T_92195 = priorityLoadRequest_3 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37651.6]
  assign _GEN_1926 = _T_92195 ? 1'h1 : loadInitiated_3; // @[AxiLoadQueue.scala 212:70:@37652.6]
  assign _GEN_1927 = initBits_3 ? 1'h0 : _GEN_1926; // @[AxiLoadQueue.scala 210:22:@37647.4]
  assign _T_92198 = priorityLoadRequest_4 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37659.6]
  assign _GEN_1928 = _T_92198 ? 1'h1 : loadInitiated_4; // @[AxiLoadQueue.scala 212:70:@37660.6]
  assign _GEN_1929 = initBits_4 ? 1'h0 : _GEN_1928; // @[AxiLoadQueue.scala 210:22:@37655.4]
  assign _T_92201 = priorityLoadRequest_5 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37667.6]
  assign _GEN_1930 = _T_92201 ? 1'h1 : loadInitiated_5; // @[AxiLoadQueue.scala 212:70:@37668.6]
  assign _GEN_1931 = initBits_5 ? 1'h0 : _GEN_1930; // @[AxiLoadQueue.scala 210:22:@37663.4]
  assign _T_92204 = priorityLoadRequest_6 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37675.6]
  assign _GEN_1932 = _T_92204 ? 1'h1 : loadInitiated_6; // @[AxiLoadQueue.scala 212:70:@37676.6]
  assign _GEN_1933 = initBits_6 ? 1'h0 : _GEN_1932; // @[AxiLoadQueue.scala 210:22:@37671.4]
  assign _T_92207 = priorityLoadRequest_7 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37683.6]
  assign _GEN_1934 = _T_92207 ? 1'h1 : loadInitiated_7; // @[AxiLoadQueue.scala 212:70:@37684.6]
  assign _GEN_1935 = initBits_7 ? 1'h0 : _GEN_1934; // @[AxiLoadQueue.scala 210:22:@37679.4]
  assign _T_92210 = priorityLoadRequest_8 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37691.6]
  assign _GEN_1936 = _T_92210 ? 1'h1 : loadInitiated_8; // @[AxiLoadQueue.scala 212:70:@37692.6]
  assign _GEN_1937 = initBits_8 ? 1'h0 : _GEN_1936; // @[AxiLoadQueue.scala 210:22:@37687.4]
  assign _T_92213 = priorityLoadRequest_9 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37699.6]
  assign _GEN_1938 = _T_92213 ? 1'h1 : loadInitiated_9; // @[AxiLoadQueue.scala 212:70:@37700.6]
  assign _GEN_1939 = initBits_9 ? 1'h0 : _GEN_1938; // @[AxiLoadQueue.scala 210:22:@37695.4]
  assign _T_92216 = priorityLoadRequest_10 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37707.6]
  assign _GEN_1940 = _T_92216 ? 1'h1 : loadInitiated_10; // @[AxiLoadQueue.scala 212:70:@37708.6]
  assign _GEN_1941 = initBits_10 ? 1'h0 : _GEN_1940; // @[AxiLoadQueue.scala 210:22:@37703.4]
  assign _T_92219 = priorityLoadRequest_11 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37715.6]
  assign _GEN_1942 = _T_92219 ? 1'h1 : loadInitiated_11; // @[AxiLoadQueue.scala 212:70:@37716.6]
  assign _GEN_1943 = initBits_11 ? 1'h0 : _GEN_1942; // @[AxiLoadQueue.scala 210:22:@37711.4]
  assign _T_92222 = priorityLoadRequest_12 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37723.6]
  assign _GEN_1944 = _T_92222 ? 1'h1 : loadInitiated_12; // @[AxiLoadQueue.scala 212:70:@37724.6]
  assign _GEN_1945 = initBits_12 ? 1'h0 : _GEN_1944; // @[AxiLoadQueue.scala 210:22:@37719.4]
  assign _T_92225 = priorityLoadRequest_13 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37731.6]
  assign _GEN_1946 = _T_92225 ? 1'h1 : loadInitiated_13; // @[AxiLoadQueue.scala 212:70:@37732.6]
  assign _GEN_1947 = initBits_13 ? 1'h0 : _GEN_1946; // @[AxiLoadQueue.scala 210:22:@37727.4]
  assign _T_92228 = priorityLoadRequest_14 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37739.6]
  assign _GEN_1948 = _T_92228 ? 1'h1 : loadInitiated_14; // @[AxiLoadQueue.scala 212:70:@37740.6]
  assign _GEN_1949 = initBits_14 ? 1'h0 : _GEN_1948; // @[AxiLoadQueue.scala 210:22:@37735.4]
  assign _T_92231 = priorityLoadRequest_15 & io_loadQIdxForAddrOut_ready; // @[AxiLoadQueue.scala 212:39:@37747.6]
  assign _GEN_1950 = _T_92231 ? 1'h1 : loadInitiated_15; // @[AxiLoadQueue.scala 212:70:@37748.6]
  assign _GEN_1951 = initBits_15 ? 1'h0 : _GEN_1950; // @[AxiLoadQueue.scala 210:22:@37743.4]
  assign _T_92249 = priorityLoadRequest_14 ? 4'he : 4'hf; // @[Mux.scala 31:69:@37751.4]
  assign _T_92250 = priorityLoadRequest_13 ? 4'hd : _T_92249; // @[Mux.scala 31:69:@37752.4]
  assign _T_92251 = priorityLoadRequest_12 ? 4'hc : _T_92250; // @[Mux.scala 31:69:@37753.4]
  assign _T_92252 = priorityLoadRequest_11 ? 4'hb : _T_92251; // @[Mux.scala 31:69:@37754.4]
  assign _T_92253 = priorityLoadRequest_10 ? 4'ha : _T_92252; // @[Mux.scala 31:69:@37755.4]
  assign _T_92254 = priorityLoadRequest_9 ? 4'h9 : _T_92253; // @[Mux.scala 31:69:@37756.4]
  assign _T_92255 = priorityLoadRequest_8 ? 4'h8 : _T_92254; // @[Mux.scala 31:69:@37757.4]
  assign _T_92256 = priorityLoadRequest_7 ? 4'h7 : _T_92255; // @[Mux.scala 31:69:@37758.4]
  assign _T_92257 = priorityLoadRequest_6 ? 4'h6 : _T_92256; // @[Mux.scala 31:69:@37759.4]
  assign _T_92258 = priorityLoadRequest_5 ? 4'h5 : _T_92257; // @[Mux.scala 31:69:@37760.4]
  assign _T_92259 = priorityLoadRequest_4 ? 4'h4 : _T_92258; // @[Mux.scala 31:69:@37761.4]
  assign _T_92260 = priorityLoadRequest_3 ? 4'h3 : _T_92259; // @[Mux.scala 31:69:@37762.4]
  assign _T_92261 = priorityLoadRequest_2 ? 4'h2 : _T_92260; // @[Mux.scala 31:69:@37763.4]
  assign _T_92262 = priorityLoadRequest_1 ? 4'h1 : _T_92261; // @[Mux.scala 31:69:@37764.4]
  assign _T_92263 = priorityLoadRequest_0 ? 4'h0 : _T_92262; // @[Mux.scala 31:69:@37765.4]
  assign _T_92266 = priorityLoadRequest_0 | priorityLoadRequest_1; // @[AxiLoadQueue.scala 222:60:@37768.4]
  assign _T_92267 = _T_92266 | priorityLoadRequest_2; // @[AxiLoadQueue.scala 222:60:@37769.4]
  assign _T_92268 = _T_92267 | priorityLoadRequest_3; // @[AxiLoadQueue.scala 222:60:@37770.4]
  assign _T_92269 = _T_92268 | priorityLoadRequest_4; // @[AxiLoadQueue.scala 222:60:@37771.4]
  assign _T_92270 = _T_92269 | priorityLoadRequest_5; // @[AxiLoadQueue.scala 222:60:@37772.4]
  assign _T_92271 = _T_92270 | priorityLoadRequest_6; // @[AxiLoadQueue.scala 222:60:@37773.4]
  assign _T_92272 = _T_92271 | priorityLoadRequest_7; // @[AxiLoadQueue.scala 222:60:@37774.4]
  assign _T_92273 = _T_92272 | priorityLoadRequest_8; // @[AxiLoadQueue.scala 222:60:@37775.4]
  assign _T_92274 = _T_92273 | priorityLoadRequest_9; // @[AxiLoadQueue.scala 222:60:@37776.4]
  assign _T_92275 = _T_92274 | priorityLoadRequest_10; // @[AxiLoadQueue.scala 222:60:@37777.4]
  assign _T_92276 = _T_92275 | priorityLoadRequest_11; // @[AxiLoadQueue.scala 222:60:@37778.4]
  assign _T_92277 = _T_92276 | priorityLoadRequest_12; // @[AxiLoadQueue.scala 222:60:@37779.4]
  assign _T_92278 = _T_92277 | priorityLoadRequest_13; // @[AxiLoadQueue.scala 222:60:@37780.4]
  assign _T_92279 = _T_92278 | priorityLoadRequest_14; // @[AxiLoadQueue.scala 222:60:@37781.4]
  assign _GEN_1953 = 4'h1 == _T_92263 ? addrQ_1 : addrQ_0; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1954 = 4'h2 == _T_92263 ? addrQ_2 : _GEN_1953; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1955 = 4'h3 == _T_92263 ? addrQ_3 : _GEN_1954; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1956 = 4'h4 == _T_92263 ? addrQ_4 : _GEN_1955; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1957 = 4'h5 == _T_92263 ? addrQ_5 : _GEN_1956; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1958 = 4'h6 == _T_92263 ? addrQ_6 : _GEN_1957; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1959 = 4'h7 == _T_92263 ? addrQ_7 : _GEN_1958; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1960 = 4'h8 == _T_92263 ? addrQ_8 : _GEN_1959; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1961 = 4'h9 == _T_92263 ? addrQ_9 : _GEN_1960; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1962 = 4'ha == _T_92263 ? addrQ_10 : _GEN_1961; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1963 = 4'hb == _T_92263 ? addrQ_11 : _GEN_1962; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1964 = 4'hc == _T_92263 ? addrQ_12 : _GEN_1963; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1965 = 4'hd == _T_92263 ? addrQ_13 : _GEN_1964; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _GEN_1966 = 4'he == _T_92263 ? addrQ_14 : _GEN_1965; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign _T_92405 = {storeAddrNotKnownFlagsPReg_0_7,storeAddrNotKnownFlagsPReg_0_6,storeAddrNotKnownFlagsPReg_0_5,storeAddrNotKnownFlagsPReg_0_4,storeAddrNotKnownFlagsPReg_0_3,storeAddrNotKnownFlagsPReg_0_2,storeAddrNotKnownFlagsPReg_0_1,storeAddrNotKnownFlagsPReg_0_0}; // @[AxiLoadQueue.scala 251:58:@37965.8]
  assign _T_92413 = {storeAddrNotKnownFlagsPReg_0_15,storeAddrNotKnownFlagsPReg_0_14,storeAddrNotKnownFlagsPReg_0_13,storeAddrNotKnownFlagsPReg_0_12,storeAddrNotKnownFlagsPReg_0_11,storeAddrNotKnownFlagsPReg_0_10,storeAddrNotKnownFlagsPReg_0_9,storeAddrNotKnownFlagsPReg_0_8,_T_92405}; // @[AxiLoadQueue.scala 251:58:@37973.8]
  assign _T_92420 = {lastConflict_0_7,lastConflict_0_6,lastConflict_0_5,lastConflict_0_4,lastConflict_0_3,lastConflict_0_2,lastConflict_0_1,lastConflict_0_0}; // @[AxiLoadQueue.scala 251:96:@37980.8]
  assign _T_92428 = {lastConflict_0_15,lastConflict_0_14,lastConflict_0_13,lastConflict_0_12,lastConflict_0_11,lastConflict_0_10,lastConflict_0_9,lastConflict_0_8,_T_92420}; // @[AxiLoadQueue.scala 251:96:@37988.8]
  assign _T_92429 = _T_92413 < _T_92428; // @[AxiLoadQueue.scala 251:61:@37989.8]
  assign _T_92430 = canBypass_0 & _T_92429; // @[AxiLoadQueue.scala 250:64:@37990.8]
  assign _GEN_2001 = _T_92359 ? _T_92430 : 1'h0; // @[AxiLoadQueue.scala 243:104:@37922.6]
  assign bypassRequest_0 = _T_92351 ? _GEN_2001 : 1'h0; // @[AxiLoadQueue.scala 242:71:@37916.4]
  assign _GEN_1968 = bypassRequest_0 ? 1'h1 : bypassInitiated_0; // @[AxiLoadQueue.scala 230:34:@37804.6]
  assign _GEN_1969 = initBits_0 ? 1'h0 : _GEN_1968; // @[AxiLoadQueue.scala 228:23:@37800.4]
  assign _T_92489 = {storeAddrNotKnownFlagsPReg_1_7,storeAddrNotKnownFlagsPReg_1_6,storeAddrNotKnownFlagsPReg_1_5,storeAddrNotKnownFlagsPReg_1_4,storeAddrNotKnownFlagsPReg_1_3,storeAddrNotKnownFlagsPReg_1_2,storeAddrNotKnownFlagsPReg_1_1,storeAddrNotKnownFlagsPReg_1_0}; // @[AxiLoadQueue.scala 251:58:@38047.8]
  assign _T_92497 = {storeAddrNotKnownFlagsPReg_1_15,storeAddrNotKnownFlagsPReg_1_14,storeAddrNotKnownFlagsPReg_1_13,storeAddrNotKnownFlagsPReg_1_12,storeAddrNotKnownFlagsPReg_1_11,storeAddrNotKnownFlagsPReg_1_10,storeAddrNotKnownFlagsPReg_1_9,storeAddrNotKnownFlagsPReg_1_8,_T_92489}; // @[AxiLoadQueue.scala 251:58:@38055.8]
  assign _T_92504 = {lastConflict_1_7,lastConflict_1_6,lastConflict_1_5,lastConflict_1_4,lastConflict_1_3,lastConflict_1_2,lastConflict_1_1,lastConflict_1_0}; // @[AxiLoadQueue.scala 251:96:@38062.8]
  assign _T_92512 = {lastConflict_1_15,lastConflict_1_14,lastConflict_1_13,lastConflict_1_12,lastConflict_1_11,lastConflict_1_10,lastConflict_1_9,lastConflict_1_8,_T_92504}; // @[AxiLoadQueue.scala 251:96:@38070.8]
  assign _T_92513 = _T_92497 < _T_92512; // @[AxiLoadQueue.scala 251:61:@38071.8]
  assign _T_92514 = canBypass_1 & _T_92513; // @[AxiLoadQueue.scala 250:64:@38072.8]
  assign _GEN_2005 = _T_92443 ? _T_92514 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38004.6]
  assign bypassRequest_1 = _T_92435 ? _GEN_2005 : 1'h0; // @[AxiLoadQueue.scala 242:71:@37998.4]
  assign _GEN_1970 = bypassRequest_1 ? 1'h1 : bypassInitiated_1; // @[AxiLoadQueue.scala 230:34:@37811.6]
  assign _GEN_1971 = initBits_1 ? 1'h0 : _GEN_1970; // @[AxiLoadQueue.scala 228:23:@37807.4]
  assign _T_92573 = {storeAddrNotKnownFlagsPReg_2_7,storeAddrNotKnownFlagsPReg_2_6,storeAddrNotKnownFlagsPReg_2_5,storeAddrNotKnownFlagsPReg_2_4,storeAddrNotKnownFlagsPReg_2_3,storeAddrNotKnownFlagsPReg_2_2,storeAddrNotKnownFlagsPReg_2_1,storeAddrNotKnownFlagsPReg_2_0}; // @[AxiLoadQueue.scala 251:58:@38129.8]
  assign _T_92581 = {storeAddrNotKnownFlagsPReg_2_15,storeAddrNotKnownFlagsPReg_2_14,storeAddrNotKnownFlagsPReg_2_13,storeAddrNotKnownFlagsPReg_2_12,storeAddrNotKnownFlagsPReg_2_11,storeAddrNotKnownFlagsPReg_2_10,storeAddrNotKnownFlagsPReg_2_9,storeAddrNotKnownFlagsPReg_2_8,_T_92573}; // @[AxiLoadQueue.scala 251:58:@38137.8]
  assign _T_92588 = {lastConflict_2_7,lastConflict_2_6,lastConflict_2_5,lastConflict_2_4,lastConflict_2_3,lastConflict_2_2,lastConflict_2_1,lastConflict_2_0}; // @[AxiLoadQueue.scala 251:96:@38144.8]
  assign _T_92596 = {lastConflict_2_15,lastConflict_2_14,lastConflict_2_13,lastConflict_2_12,lastConflict_2_11,lastConflict_2_10,lastConflict_2_9,lastConflict_2_8,_T_92588}; // @[AxiLoadQueue.scala 251:96:@38152.8]
  assign _T_92597 = _T_92581 < _T_92596; // @[AxiLoadQueue.scala 251:61:@38153.8]
  assign _T_92598 = canBypass_2 & _T_92597; // @[AxiLoadQueue.scala 250:64:@38154.8]
  assign _GEN_2009 = _T_92527 ? _T_92598 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38086.6]
  assign bypassRequest_2 = _T_92519 ? _GEN_2009 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38080.4]
  assign _GEN_1972 = bypassRequest_2 ? 1'h1 : bypassInitiated_2; // @[AxiLoadQueue.scala 230:34:@37818.6]
  assign _GEN_1973 = initBits_2 ? 1'h0 : _GEN_1972; // @[AxiLoadQueue.scala 228:23:@37814.4]
  assign _T_92657 = {storeAddrNotKnownFlagsPReg_3_7,storeAddrNotKnownFlagsPReg_3_6,storeAddrNotKnownFlagsPReg_3_5,storeAddrNotKnownFlagsPReg_3_4,storeAddrNotKnownFlagsPReg_3_3,storeAddrNotKnownFlagsPReg_3_2,storeAddrNotKnownFlagsPReg_3_1,storeAddrNotKnownFlagsPReg_3_0}; // @[AxiLoadQueue.scala 251:58:@38211.8]
  assign _T_92665 = {storeAddrNotKnownFlagsPReg_3_15,storeAddrNotKnownFlagsPReg_3_14,storeAddrNotKnownFlagsPReg_3_13,storeAddrNotKnownFlagsPReg_3_12,storeAddrNotKnownFlagsPReg_3_11,storeAddrNotKnownFlagsPReg_3_10,storeAddrNotKnownFlagsPReg_3_9,storeAddrNotKnownFlagsPReg_3_8,_T_92657}; // @[AxiLoadQueue.scala 251:58:@38219.8]
  assign _T_92672 = {lastConflict_3_7,lastConflict_3_6,lastConflict_3_5,lastConflict_3_4,lastConflict_3_3,lastConflict_3_2,lastConflict_3_1,lastConflict_3_0}; // @[AxiLoadQueue.scala 251:96:@38226.8]
  assign _T_92680 = {lastConflict_3_15,lastConflict_3_14,lastConflict_3_13,lastConflict_3_12,lastConflict_3_11,lastConflict_3_10,lastConflict_3_9,lastConflict_3_8,_T_92672}; // @[AxiLoadQueue.scala 251:96:@38234.8]
  assign _T_92681 = _T_92665 < _T_92680; // @[AxiLoadQueue.scala 251:61:@38235.8]
  assign _T_92682 = canBypass_3 & _T_92681; // @[AxiLoadQueue.scala 250:64:@38236.8]
  assign _GEN_2013 = _T_92611 ? _T_92682 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38168.6]
  assign bypassRequest_3 = _T_92603 ? _GEN_2013 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38162.4]
  assign _GEN_1974 = bypassRequest_3 ? 1'h1 : bypassInitiated_3; // @[AxiLoadQueue.scala 230:34:@37825.6]
  assign _GEN_1975 = initBits_3 ? 1'h0 : _GEN_1974; // @[AxiLoadQueue.scala 228:23:@37821.4]
  assign _T_92741 = {storeAddrNotKnownFlagsPReg_4_7,storeAddrNotKnownFlagsPReg_4_6,storeAddrNotKnownFlagsPReg_4_5,storeAddrNotKnownFlagsPReg_4_4,storeAddrNotKnownFlagsPReg_4_3,storeAddrNotKnownFlagsPReg_4_2,storeAddrNotKnownFlagsPReg_4_1,storeAddrNotKnownFlagsPReg_4_0}; // @[AxiLoadQueue.scala 251:58:@38293.8]
  assign _T_92749 = {storeAddrNotKnownFlagsPReg_4_15,storeAddrNotKnownFlagsPReg_4_14,storeAddrNotKnownFlagsPReg_4_13,storeAddrNotKnownFlagsPReg_4_12,storeAddrNotKnownFlagsPReg_4_11,storeAddrNotKnownFlagsPReg_4_10,storeAddrNotKnownFlagsPReg_4_9,storeAddrNotKnownFlagsPReg_4_8,_T_92741}; // @[AxiLoadQueue.scala 251:58:@38301.8]
  assign _T_92756 = {lastConflict_4_7,lastConflict_4_6,lastConflict_4_5,lastConflict_4_4,lastConflict_4_3,lastConflict_4_2,lastConflict_4_1,lastConflict_4_0}; // @[AxiLoadQueue.scala 251:96:@38308.8]
  assign _T_92764 = {lastConflict_4_15,lastConflict_4_14,lastConflict_4_13,lastConflict_4_12,lastConflict_4_11,lastConflict_4_10,lastConflict_4_9,lastConflict_4_8,_T_92756}; // @[AxiLoadQueue.scala 251:96:@38316.8]
  assign _T_92765 = _T_92749 < _T_92764; // @[AxiLoadQueue.scala 251:61:@38317.8]
  assign _T_92766 = canBypass_4 & _T_92765; // @[AxiLoadQueue.scala 250:64:@38318.8]
  assign _GEN_2017 = _T_92695 ? _T_92766 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38250.6]
  assign bypassRequest_4 = _T_92687 ? _GEN_2017 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38244.4]
  assign _GEN_1976 = bypassRequest_4 ? 1'h1 : bypassInitiated_4; // @[AxiLoadQueue.scala 230:34:@37832.6]
  assign _GEN_1977 = initBits_4 ? 1'h0 : _GEN_1976; // @[AxiLoadQueue.scala 228:23:@37828.4]
  assign _T_92825 = {storeAddrNotKnownFlagsPReg_5_7,storeAddrNotKnownFlagsPReg_5_6,storeAddrNotKnownFlagsPReg_5_5,storeAddrNotKnownFlagsPReg_5_4,storeAddrNotKnownFlagsPReg_5_3,storeAddrNotKnownFlagsPReg_5_2,storeAddrNotKnownFlagsPReg_5_1,storeAddrNotKnownFlagsPReg_5_0}; // @[AxiLoadQueue.scala 251:58:@38375.8]
  assign _T_92833 = {storeAddrNotKnownFlagsPReg_5_15,storeAddrNotKnownFlagsPReg_5_14,storeAddrNotKnownFlagsPReg_5_13,storeAddrNotKnownFlagsPReg_5_12,storeAddrNotKnownFlagsPReg_5_11,storeAddrNotKnownFlagsPReg_5_10,storeAddrNotKnownFlagsPReg_5_9,storeAddrNotKnownFlagsPReg_5_8,_T_92825}; // @[AxiLoadQueue.scala 251:58:@38383.8]
  assign _T_92840 = {lastConflict_5_7,lastConflict_5_6,lastConflict_5_5,lastConflict_5_4,lastConflict_5_3,lastConflict_5_2,lastConflict_5_1,lastConflict_5_0}; // @[AxiLoadQueue.scala 251:96:@38390.8]
  assign _T_92848 = {lastConflict_5_15,lastConflict_5_14,lastConflict_5_13,lastConflict_5_12,lastConflict_5_11,lastConflict_5_10,lastConflict_5_9,lastConflict_5_8,_T_92840}; // @[AxiLoadQueue.scala 251:96:@38398.8]
  assign _T_92849 = _T_92833 < _T_92848; // @[AxiLoadQueue.scala 251:61:@38399.8]
  assign _T_92850 = canBypass_5 & _T_92849; // @[AxiLoadQueue.scala 250:64:@38400.8]
  assign _GEN_2021 = _T_92779 ? _T_92850 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38332.6]
  assign bypassRequest_5 = _T_92771 ? _GEN_2021 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38326.4]
  assign _GEN_1978 = bypassRequest_5 ? 1'h1 : bypassInitiated_5; // @[AxiLoadQueue.scala 230:34:@37839.6]
  assign _GEN_1979 = initBits_5 ? 1'h0 : _GEN_1978; // @[AxiLoadQueue.scala 228:23:@37835.4]
  assign _T_92909 = {storeAddrNotKnownFlagsPReg_6_7,storeAddrNotKnownFlagsPReg_6_6,storeAddrNotKnownFlagsPReg_6_5,storeAddrNotKnownFlagsPReg_6_4,storeAddrNotKnownFlagsPReg_6_3,storeAddrNotKnownFlagsPReg_6_2,storeAddrNotKnownFlagsPReg_6_1,storeAddrNotKnownFlagsPReg_6_0}; // @[AxiLoadQueue.scala 251:58:@38457.8]
  assign _T_92917 = {storeAddrNotKnownFlagsPReg_6_15,storeAddrNotKnownFlagsPReg_6_14,storeAddrNotKnownFlagsPReg_6_13,storeAddrNotKnownFlagsPReg_6_12,storeAddrNotKnownFlagsPReg_6_11,storeAddrNotKnownFlagsPReg_6_10,storeAddrNotKnownFlagsPReg_6_9,storeAddrNotKnownFlagsPReg_6_8,_T_92909}; // @[AxiLoadQueue.scala 251:58:@38465.8]
  assign _T_92924 = {lastConflict_6_7,lastConflict_6_6,lastConflict_6_5,lastConflict_6_4,lastConflict_6_3,lastConflict_6_2,lastConflict_6_1,lastConflict_6_0}; // @[AxiLoadQueue.scala 251:96:@38472.8]
  assign _T_92932 = {lastConflict_6_15,lastConflict_6_14,lastConflict_6_13,lastConflict_6_12,lastConflict_6_11,lastConflict_6_10,lastConflict_6_9,lastConflict_6_8,_T_92924}; // @[AxiLoadQueue.scala 251:96:@38480.8]
  assign _T_92933 = _T_92917 < _T_92932; // @[AxiLoadQueue.scala 251:61:@38481.8]
  assign _T_92934 = canBypass_6 & _T_92933; // @[AxiLoadQueue.scala 250:64:@38482.8]
  assign _GEN_2025 = _T_92863 ? _T_92934 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38414.6]
  assign bypassRequest_6 = _T_92855 ? _GEN_2025 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38408.4]
  assign _GEN_1980 = bypassRequest_6 ? 1'h1 : bypassInitiated_6; // @[AxiLoadQueue.scala 230:34:@37846.6]
  assign _GEN_1981 = initBits_6 ? 1'h0 : _GEN_1980; // @[AxiLoadQueue.scala 228:23:@37842.4]
  assign _T_92993 = {storeAddrNotKnownFlagsPReg_7_7,storeAddrNotKnownFlagsPReg_7_6,storeAddrNotKnownFlagsPReg_7_5,storeAddrNotKnownFlagsPReg_7_4,storeAddrNotKnownFlagsPReg_7_3,storeAddrNotKnownFlagsPReg_7_2,storeAddrNotKnownFlagsPReg_7_1,storeAddrNotKnownFlagsPReg_7_0}; // @[AxiLoadQueue.scala 251:58:@38539.8]
  assign _T_93001 = {storeAddrNotKnownFlagsPReg_7_15,storeAddrNotKnownFlagsPReg_7_14,storeAddrNotKnownFlagsPReg_7_13,storeAddrNotKnownFlagsPReg_7_12,storeAddrNotKnownFlagsPReg_7_11,storeAddrNotKnownFlagsPReg_7_10,storeAddrNotKnownFlagsPReg_7_9,storeAddrNotKnownFlagsPReg_7_8,_T_92993}; // @[AxiLoadQueue.scala 251:58:@38547.8]
  assign _T_93008 = {lastConflict_7_7,lastConflict_7_6,lastConflict_7_5,lastConflict_7_4,lastConflict_7_3,lastConflict_7_2,lastConflict_7_1,lastConflict_7_0}; // @[AxiLoadQueue.scala 251:96:@38554.8]
  assign _T_93016 = {lastConflict_7_15,lastConflict_7_14,lastConflict_7_13,lastConflict_7_12,lastConflict_7_11,lastConflict_7_10,lastConflict_7_9,lastConflict_7_8,_T_93008}; // @[AxiLoadQueue.scala 251:96:@38562.8]
  assign _T_93017 = _T_93001 < _T_93016; // @[AxiLoadQueue.scala 251:61:@38563.8]
  assign _T_93018 = canBypass_7 & _T_93017; // @[AxiLoadQueue.scala 250:64:@38564.8]
  assign _GEN_2029 = _T_92947 ? _T_93018 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38496.6]
  assign bypassRequest_7 = _T_92939 ? _GEN_2029 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38490.4]
  assign _GEN_1982 = bypassRequest_7 ? 1'h1 : bypassInitiated_7; // @[AxiLoadQueue.scala 230:34:@37853.6]
  assign _GEN_1983 = initBits_7 ? 1'h0 : _GEN_1982; // @[AxiLoadQueue.scala 228:23:@37849.4]
  assign _T_93077 = {storeAddrNotKnownFlagsPReg_8_7,storeAddrNotKnownFlagsPReg_8_6,storeAddrNotKnownFlagsPReg_8_5,storeAddrNotKnownFlagsPReg_8_4,storeAddrNotKnownFlagsPReg_8_3,storeAddrNotKnownFlagsPReg_8_2,storeAddrNotKnownFlagsPReg_8_1,storeAddrNotKnownFlagsPReg_8_0}; // @[AxiLoadQueue.scala 251:58:@38621.8]
  assign _T_93085 = {storeAddrNotKnownFlagsPReg_8_15,storeAddrNotKnownFlagsPReg_8_14,storeAddrNotKnownFlagsPReg_8_13,storeAddrNotKnownFlagsPReg_8_12,storeAddrNotKnownFlagsPReg_8_11,storeAddrNotKnownFlagsPReg_8_10,storeAddrNotKnownFlagsPReg_8_9,storeAddrNotKnownFlagsPReg_8_8,_T_93077}; // @[AxiLoadQueue.scala 251:58:@38629.8]
  assign _T_93092 = {lastConflict_8_7,lastConflict_8_6,lastConflict_8_5,lastConflict_8_4,lastConflict_8_3,lastConflict_8_2,lastConflict_8_1,lastConflict_8_0}; // @[AxiLoadQueue.scala 251:96:@38636.8]
  assign _T_93100 = {lastConflict_8_15,lastConflict_8_14,lastConflict_8_13,lastConflict_8_12,lastConflict_8_11,lastConflict_8_10,lastConflict_8_9,lastConflict_8_8,_T_93092}; // @[AxiLoadQueue.scala 251:96:@38644.8]
  assign _T_93101 = _T_93085 < _T_93100; // @[AxiLoadQueue.scala 251:61:@38645.8]
  assign _T_93102 = canBypass_8 & _T_93101; // @[AxiLoadQueue.scala 250:64:@38646.8]
  assign _GEN_2033 = _T_93031 ? _T_93102 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38578.6]
  assign bypassRequest_8 = _T_93023 ? _GEN_2033 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38572.4]
  assign _GEN_1984 = bypassRequest_8 ? 1'h1 : bypassInitiated_8; // @[AxiLoadQueue.scala 230:34:@37860.6]
  assign _GEN_1985 = initBits_8 ? 1'h0 : _GEN_1984; // @[AxiLoadQueue.scala 228:23:@37856.4]
  assign _T_93161 = {storeAddrNotKnownFlagsPReg_9_7,storeAddrNotKnownFlagsPReg_9_6,storeAddrNotKnownFlagsPReg_9_5,storeAddrNotKnownFlagsPReg_9_4,storeAddrNotKnownFlagsPReg_9_3,storeAddrNotKnownFlagsPReg_9_2,storeAddrNotKnownFlagsPReg_9_1,storeAddrNotKnownFlagsPReg_9_0}; // @[AxiLoadQueue.scala 251:58:@38703.8]
  assign _T_93169 = {storeAddrNotKnownFlagsPReg_9_15,storeAddrNotKnownFlagsPReg_9_14,storeAddrNotKnownFlagsPReg_9_13,storeAddrNotKnownFlagsPReg_9_12,storeAddrNotKnownFlagsPReg_9_11,storeAddrNotKnownFlagsPReg_9_10,storeAddrNotKnownFlagsPReg_9_9,storeAddrNotKnownFlagsPReg_9_8,_T_93161}; // @[AxiLoadQueue.scala 251:58:@38711.8]
  assign _T_93176 = {lastConflict_9_7,lastConflict_9_6,lastConflict_9_5,lastConflict_9_4,lastConflict_9_3,lastConflict_9_2,lastConflict_9_1,lastConflict_9_0}; // @[AxiLoadQueue.scala 251:96:@38718.8]
  assign _T_93184 = {lastConflict_9_15,lastConflict_9_14,lastConflict_9_13,lastConflict_9_12,lastConflict_9_11,lastConflict_9_10,lastConflict_9_9,lastConflict_9_8,_T_93176}; // @[AxiLoadQueue.scala 251:96:@38726.8]
  assign _T_93185 = _T_93169 < _T_93184; // @[AxiLoadQueue.scala 251:61:@38727.8]
  assign _T_93186 = canBypass_9 & _T_93185; // @[AxiLoadQueue.scala 250:64:@38728.8]
  assign _GEN_2037 = _T_93115 ? _T_93186 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38660.6]
  assign bypassRequest_9 = _T_93107 ? _GEN_2037 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38654.4]
  assign _GEN_1986 = bypassRequest_9 ? 1'h1 : bypassInitiated_9; // @[AxiLoadQueue.scala 230:34:@37867.6]
  assign _GEN_1987 = initBits_9 ? 1'h0 : _GEN_1986; // @[AxiLoadQueue.scala 228:23:@37863.4]
  assign _T_93245 = {storeAddrNotKnownFlagsPReg_10_7,storeAddrNotKnownFlagsPReg_10_6,storeAddrNotKnownFlagsPReg_10_5,storeAddrNotKnownFlagsPReg_10_4,storeAddrNotKnownFlagsPReg_10_3,storeAddrNotKnownFlagsPReg_10_2,storeAddrNotKnownFlagsPReg_10_1,storeAddrNotKnownFlagsPReg_10_0}; // @[AxiLoadQueue.scala 251:58:@38785.8]
  assign _T_93253 = {storeAddrNotKnownFlagsPReg_10_15,storeAddrNotKnownFlagsPReg_10_14,storeAddrNotKnownFlagsPReg_10_13,storeAddrNotKnownFlagsPReg_10_12,storeAddrNotKnownFlagsPReg_10_11,storeAddrNotKnownFlagsPReg_10_10,storeAddrNotKnownFlagsPReg_10_9,storeAddrNotKnownFlagsPReg_10_8,_T_93245}; // @[AxiLoadQueue.scala 251:58:@38793.8]
  assign _T_93260 = {lastConflict_10_7,lastConflict_10_6,lastConflict_10_5,lastConflict_10_4,lastConflict_10_3,lastConflict_10_2,lastConflict_10_1,lastConflict_10_0}; // @[AxiLoadQueue.scala 251:96:@38800.8]
  assign _T_93268 = {lastConflict_10_15,lastConflict_10_14,lastConflict_10_13,lastConflict_10_12,lastConflict_10_11,lastConflict_10_10,lastConflict_10_9,lastConflict_10_8,_T_93260}; // @[AxiLoadQueue.scala 251:96:@38808.8]
  assign _T_93269 = _T_93253 < _T_93268; // @[AxiLoadQueue.scala 251:61:@38809.8]
  assign _T_93270 = canBypass_10 & _T_93269; // @[AxiLoadQueue.scala 250:64:@38810.8]
  assign _GEN_2041 = _T_93199 ? _T_93270 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38742.6]
  assign bypassRequest_10 = _T_93191 ? _GEN_2041 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38736.4]
  assign _GEN_1988 = bypassRequest_10 ? 1'h1 : bypassInitiated_10; // @[AxiLoadQueue.scala 230:34:@37874.6]
  assign _GEN_1989 = initBits_10 ? 1'h0 : _GEN_1988; // @[AxiLoadQueue.scala 228:23:@37870.4]
  assign _T_93329 = {storeAddrNotKnownFlagsPReg_11_7,storeAddrNotKnownFlagsPReg_11_6,storeAddrNotKnownFlagsPReg_11_5,storeAddrNotKnownFlagsPReg_11_4,storeAddrNotKnownFlagsPReg_11_3,storeAddrNotKnownFlagsPReg_11_2,storeAddrNotKnownFlagsPReg_11_1,storeAddrNotKnownFlagsPReg_11_0}; // @[AxiLoadQueue.scala 251:58:@38867.8]
  assign _T_93337 = {storeAddrNotKnownFlagsPReg_11_15,storeAddrNotKnownFlagsPReg_11_14,storeAddrNotKnownFlagsPReg_11_13,storeAddrNotKnownFlagsPReg_11_12,storeAddrNotKnownFlagsPReg_11_11,storeAddrNotKnownFlagsPReg_11_10,storeAddrNotKnownFlagsPReg_11_9,storeAddrNotKnownFlagsPReg_11_8,_T_93329}; // @[AxiLoadQueue.scala 251:58:@38875.8]
  assign _T_93344 = {lastConflict_11_7,lastConflict_11_6,lastConflict_11_5,lastConflict_11_4,lastConflict_11_3,lastConflict_11_2,lastConflict_11_1,lastConflict_11_0}; // @[AxiLoadQueue.scala 251:96:@38882.8]
  assign _T_93352 = {lastConflict_11_15,lastConflict_11_14,lastConflict_11_13,lastConflict_11_12,lastConflict_11_11,lastConflict_11_10,lastConflict_11_9,lastConflict_11_8,_T_93344}; // @[AxiLoadQueue.scala 251:96:@38890.8]
  assign _T_93353 = _T_93337 < _T_93352; // @[AxiLoadQueue.scala 251:61:@38891.8]
  assign _T_93354 = canBypass_11 & _T_93353; // @[AxiLoadQueue.scala 250:64:@38892.8]
  assign _GEN_2045 = _T_93283 ? _T_93354 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38824.6]
  assign bypassRequest_11 = _T_93275 ? _GEN_2045 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38818.4]
  assign _GEN_1990 = bypassRequest_11 ? 1'h1 : bypassInitiated_11; // @[AxiLoadQueue.scala 230:34:@37881.6]
  assign _GEN_1991 = initBits_11 ? 1'h0 : _GEN_1990; // @[AxiLoadQueue.scala 228:23:@37877.4]
  assign _T_93413 = {storeAddrNotKnownFlagsPReg_12_7,storeAddrNotKnownFlagsPReg_12_6,storeAddrNotKnownFlagsPReg_12_5,storeAddrNotKnownFlagsPReg_12_4,storeAddrNotKnownFlagsPReg_12_3,storeAddrNotKnownFlagsPReg_12_2,storeAddrNotKnownFlagsPReg_12_1,storeAddrNotKnownFlagsPReg_12_0}; // @[AxiLoadQueue.scala 251:58:@38949.8]
  assign _T_93421 = {storeAddrNotKnownFlagsPReg_12_15,storeAddrNotKnownFlagsPReg_12_14,storeAddrNotKnownFlagsPReg_12_13,storeAddrNotKnownFlagsPReg_12_12,storeAddrNotKnownFlagsPReg_12_11,storeAddrNotKnownFlagsPReg_12_10,storeAddrNotKnownFlagsPReg_12_9,storeAddrNotKnownFlagsPReg_12_8,_T_93413}; // @[AxiLoadQueue.scala 251:58:@38957.8]
  assign _T_93428 = {lastConflict_12_7,lastConflict_12_6,lastConflict_12_5,lastConflict_12_4,lastConflict_12_3,lastConflict_12_2,lastConflict_12_1,lastConflict_12_0}; // @[AxiLoadQueue.scala 251:96:@38964.8]
  assign _T_93436 = {lastConflict_12_15,lastConflict_12_14,lastConflict_12_13,lastConflict_12_12,lastConflict_12_11,lastConflict_12_10,lastConflict_12_9,lastConflict_12_8,_T_93428}; // @[AxiLoadQueue.scala 251:96:@38972.8]
  assign _T_93437 = _T_93421 < _T_93436; // @[AxiLoadQueue.scala 251:61:@38973.8]
  assign _T_93438 = canBypass_12 & _T_93437; // @[AxiLoadQueue.scala 250:64:@38974.8]
  assign _GEN_2049 = _T_93367 ? _T_93438 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38906.6]
  assign bypassRequest_12 = _T_93359 ? _GEN_2049 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38900.4]
  assign _GEN_1992 = bypassRequest_12 ? 1'h1 : bypassInitiated_12; // @[AxiLoadQueue.scala 230:34:@37888.6]
  assign _GEN_1993 = initBits_12 ? 1'h0 : _GEN_1992; // @[AxiLoadQueue.scala 228:23:@37884.4]
  assign _T_93497 = {storeAddrNotKnownFlagsPReg_13_7,storeAddrNotKnownFlagsPReg_13_6,storeAddrNotKnownFlagsPReg_13_5,storeAddrNotKnownFlagsPReg_13_4,storeAddrNotKnownFlagsPReg_13_3,storeAddrNotKnownFlagsPReg_13_2,storeAddrNotKnownFlagsPReg_13_1,storeAddrNotKnownFlagsPReg_13_0}; // @[AxiLoadQueue.scala 251:58:@39031.8]
  assign _T_93505 = {storeAddrNotKnownFlagsPReg_13_15,storeAddrNotKnownFlagsPReg_13_14,storeAddrNotKnownFlagsPReg_13_13,storeAddrNotKnownFlagsPReg_13_12,storeAddrNotKnownFlagsPReg_13_11,storeAddrNotKnownFlagsPReg_13_10,storeAddrNotKnownFlagsPReg_13_9,storeAddrNotKnownFlagsPReg_13_8,_T_93497}; // @[AxiLoadQueue.scala 251:58:@39039.8]
  assign _T_93512 = {lastConflict_13_7,lastConflict_13_6,lastConflict_13_5,lastConflict_13_4,lastConflict_13_3,lastConflict_13_2,lastConflict_13_1,lastConflict_13_0}; // @[AxiLoadQueue.scala 251:96:@39046.8]
  assign _T_93520 = {lastConflict_13_15,lastConflict_13_14,lastConflict_13_13,lastConflict_13_12,lastConflict_13_11,lastConflict_13_10,lastConflict_13_9,lastConflict_13_8,_T_93512}; // @[AxiLoadQueue.scala 251:96:@39054.8]
  assign _T_93521 = _T_93505 < _T_93520; // @[AxiLoadQueue.scala 251:61:@39055.8]
  assign _T_93522 = canBypass_13 & _T_93521; // @[AxiLoadQueue.scala 250:64:@39056.8]
  assign _GEN_2053 = _T_93451 ? _T_93522 : 1'h0; // @[AxiLoadQueue.scala 243:104:@38988.6]
  assign bypassRequest_13 = _T_93443 ? _GEN_2053 : 1'h0; // @[AxiLoadQueue.scala 242:71:@38982.4]
  assign _GEN_1994 = bypassRequest_13 ? 1'h1 : bypassInitiated_13; // @[AxiLoadQueue.scala 230:34:@37895.6]
  assign _GEN_1995 = initBits_13 ? 1'h0 : _GEN_1994; // @[AxiLoadQueue.scala 228:23:@37891.4]
  assign _T_93581 = {storeAddrNotKnownFlagsPReg_14_7,storeAddrNotKnownFlagsPReg_14_6,storeAddrNotKnownFlagsPReg_14_5,storeAddrNotKnownFlagsPReg_14_4,storeAddrNotKnownFlagsPReg_14_3,storeAddrNotKnownFlagsPReg_14_2,storeAddrNotKnownFlagsPReg_14_1,storeAddrNotKnownFlagsPReg_14_0}; // @[AxiLoadQueue.scala 251:58:@39113.8]
  assign _T_93589 = {storeAddrNotKnownFlagsPReg_14_15,storeAddrNotKnownFlagsPReg_14_14,storeAddrNotKnownFlagsPReg_14_13,storeAddrNotKnownFlagsPReg_14_12,storeAddrNotKnownFlagsPReg_14_11,storeAddrNotKnownFlagsPReg_14_10,storeAddrNotKnownFlagsPReg_14_9,storeAddrNotKnownFlagsPReg_14_8,_T_93581}; // @[AxiLoadQueue.scala 251:58:@39121.8]
  assign _T_93596 = {lastConflict_14_7,lastConflict_14_6,lastConflict_14_5,lastConflict_14_4,lastConflict_14_3,lastConflict_14_2,lastConflict_14_1,lastConflict_14_0}; // @[AxiLoadQueue.scala 251:96:@39128.8]
  assign _T_93604 = {lastConflict_14_15,lastConflict_14_14,lastConflict_14_13,lastConflict_14_12,lastConflict_14_11,lastConflict_14_10,lastConflict_14_9,lastConflict_14_8,_T_93596}; // @[AxiLoadQueue.scala 251:96:@39136.8]
  assign _T_93605 = _T_93589 < _T_93604; // @[AxiLoadQueue.scala 251:61:@39137.8]
  assign _T_93606 = canBypass_14 & _T_93605; // @[AxiLoadQueue.scala 250:64:@39138.8]
  assign _GEN_2057 = _T_93535 ? _T_93606 : 1'h0; // @[AxiLoadQueue.scala 243:104:@39070.6]
  assign bypassRequest_14 = _T_93527 ? _GEN_2057 : 1'h0; // @[AxiLoadQueue.scala 242:71:@39064.4]
  assign _GEN_1996 = bypassRequest_14 ? 1'h1 : bypassInitiated_14; // @[AxiLoadQueue.scala 230:34:@37902.6]
  assign _GEN_1997 = initBits_14 ? 1'h0 : _GEN_1996; // @[AxiLoadQueue.scala 228:23:@37898.4]
  assign _T_93665 = {storeAddrNotKnownFlagsPReg_15_7,storeAddrNotKnownFlagsPReg_15_6,storeAddrNotKnownFlagsPReg_15_5,storeAddrNotKnownFlagsPReg_15_4,storeAddrNotKnownFlagsPReg_15_3,storeAddrNotKnownFlagsPReg_15_2,storeAddrNotKnownFlagsPReg_15_1,storeAddrNotKnownFlagsPReg_15_0}; // @[AxiLoadQueue.scala 251:58:@39195.8]
  assign _T_93673 = {storeAddrNotKnownFlagsPReg_15_15,storeAddrNotKnownFlagsPReg_15_14,storeAddrNotKnownFlagsPReg_15_13,storeAddrNotKnownFlagsPReg_15_12,storeAddrNotKnownFlagsPReg_15_11,storeAddrNotKnownFlagsPReg_15_10,storeAddrNotKnownFlagsPReg_15_9,storeAddrNotKnownFlagsPReg_15_8,_T_93665}; // @[AxiLoadQueue.scala 251:58:@39203.8]
  assign _T_93680 = {lastConflict_15_7,lastConflict_15_6,lastConflict_15_5,lastConflict_15_4,lastConflict_15_3,lastConflict_15_2,lastConflict_15_1,lastConflict_15_0}; // @[AxiLoadQueue.scala 251:96:@39210.8]
  assign _T_93688 = {lastConflict_15_15,lastConflict_15_14,lastConflict_15_13,lastConflict_15_12,lastConflict_15_11,lastConflict_15_10,lastConflict_15_9,lastConflict_15_8,_T_93680}; // @[AxiLoadQueue.scala 251:96:@39218.8]
  assign _T_93689 = _T_93673 < _T_93688; // @[AxiLoadQueue.scala 251:61:@39219.8]
  assign _T_93690 = canBypass_15 & _T_93689; // @[AxiLoadQueue.scala 250:64:@39220.8]
  assign _GEN_2061 = _T_93619 ? _T_93690 : 1'h0; // @[AxiLoadQueue.scala 243:104:@39152.6]
  assign bypassRequest_15 = _T_93611 ? _GEN_2061 : 1'h0; // @[AxiLoadQueue.scala 242:71:@39146.4]
  assign _GEN_1998 = bypassRequest_15 ? 1'h1 : bypassInitiated_15; // @[AxiLoadQueue.scala 230:34:@37909.6]
  assign _GEN_1999 = initBits_15 ? 1'h0 : _GEN_1998; // @[AxiLoadQueue.scala 228:23:@37905.4]
  assign _T_93693 = io_loadQIdxForDataIn == 32'h0; // @[AxiLoadQueue.scala 262:69:@39228.6]
  assign _T_93694 = io_loadQIdxForDataInValid & _T_93693; // @[AxiLoadQueue.scala 262:45:@39229.6]
  assign _T_93695 = _T_93694 | bypassRequest_0; // @[AxiLoadQueue.scala 262:78:@39230.6]
  assign _GEN_2064 = _T_93695 ? 1'h1 : dataKnown_0; // @[AxiLoadQueue.scala 262:99:@39231.6]
  assign _GEN_2065 = initBits_0 ? 1'h0 : _GEN_2064; // @[AxiLoadQueue.scala 260:25:@39224.4]
  assign _T_93699 = io_loadQIdxForDataIn == 32'h1; // @[AxiLoadQueue.scala 262:69:@39238.6]
  assign _T_93700 = io_loadQIdxForDataInValid & _T_93699; // @[AxiLoadQueue.scala 262:45:@39239.6]
  assign _T_93701 = _T_93700 | bypassRequest_1; // @[AxiLoadQueue.scala 262:78:@39240.6]
  assign _GEN_2066 = _T_93701 ? 1'h1 : dataKnown_1; // @[AxiLoadQueue.scala 262:99:@39241.6]
  assign _GEN_2067 = initBits_1 ? 1'h0 : _GEN_2066; // @[AxiLoadQueue.scala 260:25:@39234.4]
  assign _T_93705 = io_loadQIdxForDataIn == 32'h2; // @[AxiLoadQueue.scala 262:69:@39248.6]
  assign _T_93706 = io_loadQIdxForDataInValid & _T_93705; // @[AxiLoadQueue.scala 262:45:@39249.6]
  assign _T_93707 = _T_93706 | bypassRequest_2; // @[AxiLoadQueue.scala 262:78:@39250.6]
  assign _GEN_2068 = _T_93707 ? 1'h1 : dataKnown_2; // @[AxiLoadQueue.scala 262:99:@39251.6]
  assign _GEN_2069 = initBits_2 ? 1'h0 : _GEN_2068; // @[AxiLoadQueue.scala 260:25:@39244.4]
  assign _T_93711 = io_loadQIdxForDataIn == 32'h3; // @[AxiLoadQueue.scala 262:69:@39258.6]
  assign _T_93712 = io_loadQIdxForDataInValid & _T_93711; // @[AxiLoadQueue.scala 262:45:@39259.6]
  assign _T_93713 = _T_93712 | bypassRequest_3; // @[AxiLoadQueue.scala 262:78:@39260.6]
  assign _GEN_2070 = _T_93713 ? 1'h1 : dataKnown_3; // @[AxiLoadQueue.scala 262:99:@39261.6]
  assign _GEN_2071 = initBits_3 ? 1'h0 : _GEN_2070; // @[AxiLoadQueue.scala 260:25:@39254.4]
  assign _T_93717 = io_loadQIdxForDataIn == 32'h4; // @[AxiLoadQueue.scala 262:69:@39268.6]
  assign _T_93718 = io_loadQIdxForDataInValid & _T_93717; // @[AxiLoadQueue.scala 262:45:@39269.6]
  assign _T_93719 = _T_93718 | bypassRequest_4; // @[AxiLoadQueue.scala 262:78:@39270.6]
  assign _GEN_2072 = _T_93719 ? 1'h1 : dataKnown_4; // @[AxiLoadQueue.scala 262:99:@39271.6]
  assign _GEN_2073 = initBits_4 ? 1'h0 : _GEN_2072; // @[AxiLoadQueue.scala 260:25:@39264.4]
  assign _T_93723 = io_loadQIdxForDataIn == 32'h5; // @[AxiLoadQueue.scala 262:69:@39278.6]
  assign _T_93724 = io_loadQIdxForDataInValid & _T_93723; // @[AxiLoadQueue.scala 262:45:@39279.6]
  assign _T_93725 = _T_93724 | bypassRequest_5; // @[AxiLoadQueue.scala 262:78:@39280.6]
  assign _GEN_2074 = _T_93725 ? 1'h1 : dataKnown_5; // @[AxiLoadQueue.scala 262:99:@39281.6]
  assign _GEN_2075 = initBits_5 ? 1'h0 : _GEN_2074; // @[AxiLoadQueue.scala 260:25:@39274.4]
  assign _T_93729 = io_loadQIdxForDataIn == 32'h6; // @[AxiLoadQueue.scala 262:69:@39288.6]
  assign _T_93730 = io_loadQIdxForDataInValid & _T_93729; // @[AxiLoadQueue.scala 262:45:@39289.6]
  assign _T_93731 = _T_93730 | bypassRequest_6; // @[AxiLoadQueue.scala 262:78:@39290.6]
  assign _GEN_2076 = _T_93731 ? 1'h1 : dataKnown_6; // @[AxiLoadQueue.scala 262:99:@39291.6]
  assign _GEN_2077 = initBits_6 ? 1'h0 : _GEN_2076; // @[AxiLoadQueue.scala 260:25:@39284.4]
  assign _T_93735 = io_loadQIdxForDataIn == 32'h7; // @[AxiLoadQueue.scala 262:69:@39298.6]
  assign _T_93736 = io_loadQIdxForDataInValid & _T_93735; // @[AxiLoadQueue.scala 262:45:@39299.6]
  assign _T_93737 = _T_93736 | bypassRequest_7; // @[AxiLoadQueue.scala 262:78:@39300.6]
  assign _GEN_2078 = _T_93737 ? 1'h1 : dataKnown_7; // @[AxiLoadQueue.scala 262:99:@39301.6]
  assign _GEN_2079 = initBits_7 ? 1'h0 : _GEN_2078; // @[AxiLoadQueue.scala 260:25:@39294.4]
  assign _T_93741 = io_loadQIdxForDataIn == 32'h8; // @[AxiLoadQueue.scala 262:69:@39308.6]
  assign _T_93742 = io_loadQIdxForDataInValid & _T_93741; // @[AxiLoadQueue.scala 262:45:@39309.6]
  assign _T_93743 = _T_93742 | bypassRequest_8; // @[AxiLoadQueue.scala 262:78:@39310.6]
  assign _GEN_2080 = _T_93743 ? 1'h1 : dataKnown_8; // @[AxiLoadQueue.scala 262:99:@39311.6]
  assign _GEN_2081 = initBits_8 ? 1'h0 : _GEN_2080; // @[AxiLoadQueue.scala 260:25:@39304.4]
  assign _T_93747 = io_loadQIdxForDataIn == 32'h9; // @[AxiLoadQueue.scala 262:69:@39318.6]
  assign _T_93748 = io_loadQIdxForDataInValid & _T_93747; // @[AxiLoadQueue.scala 262:45:@39319.6]
  assign _T_93749 = _T_93748 | bypassRequest_9; // @[AxiLoadQueue.scala 262:78:@39320.6]
  assign _GEN_2082 = _T_93749 ? 1'h1 : dataKnown_9; // @[AxiLoadQueue.scala 262:99:@39321.6]
  assign _GEN_2083 = initBits_9 ? 1'h0 : _GEN_2082; // @[AxiLoadQueue.scala 260:25:@39314.4]
  assign _T_93753 = io_loadQIdxForDataIn == 32'ha; // @[AxiLoadQueue.scala 262:69:@39328.6]
  assign _T_93754 = io_loadQIdxForDataInValid & _T_93753; // @[AxiLoadQueue.scala 262:45:@39329.6]
  assign _T_93755 = _T_93754 | bypassRequest_10; // @[AxiLoadQueue.scala 262:78:@39330.6]
  assign _GEN_2084 = _T_93755 ? 1'h1 : dataKnown_10; // @[AxiLoadQueue.scala 262:99:@39331.6]
  assign _GEN_2085 = initBits_10 ? 1'h0 : _GEN_2084; // @[AxiLoadQueue.scala 260:25:@39324.4]
  assign _T_93759 = io_loadQIdxForDataIn == 32'hb; // @[AxiLoadQueue.scala 262:69:@39338.6]
  assign _T_93760 = io_loadQIdxForDataInValid & _T_93759; // @[AxiLoadQueue.scala 262:45:@39339.6]
  assign _T_93761 = _T_93760 | bypassRequest_11; // @[AxiLoadQueue.scala 262:78:@39340.6]
  assign _GEN_2086 = _T_93761 ? 1'h1 : dataKnown_11; // @[AxiLoadQueue.scala 262:99:@39341.6]
  assign _GEN_2087 = initBits_11 ? 1'h0 : _GEN_2086; // @[AxiLoadQueue.scala 260:25:@39334.4]
  assign _T_93765 = io_loadQIdxForDataIn == 32'hc; // @[AxiLoadQueue.scala 262:69:@39348.6]
  assign _T_93766 = io_loadQIdxForDataInValid & _T_93765; // @[AxiLoadQueue.scala 262:45:@39349.6]
  assign _T_93767 = _T_93766 | bypassRequest_12; // @[AxiLoadQueue.scala 262:78:@39350.6]
  assign _GEN_2088 = _T_93767 ? 1'h1 : dataKnown_12; // @[AxiLoadQueue.scala 262:99:@39351.6]
  assign _GEN_2089 = initBits_12 ? 1'h0 : _GEN_2088; // @[AxiLoadQueue.scala 260:25:@39344.4]
  assign _T_93771 = io_loadQIdxForDataIn == 32'hd; // @[AxiLoadQueue.scala 262:69:@39358.6]
  assign _T_93772 = io_loadQIdxForDataInValid & _T_93771; // @[AxiLoadQueue.scala 262:45:@39359.6]
  assign _T_93773 = _T_93772 | bypassRequest_13; // @[AxiLoadQueue.scala 262:78:@39360.6]
  assign _GEN_2090 = _T_93773 ? 1'h1 : dataKnown_13; // @[AxiLoadQueue.scala 262:99:@39361.6]
  assign _GEN_2091 = initBits_13 ? 1'h0 : _GEN_2090; // @[AxiLoadQueue.scala 260:25:@39354.4]
  assign _T_93777 = io_loadQIdxForDataIn == 32'he; // @[AxiLoadQueue.scala 262:69:@39368.6]
  assign _T_93778 = io_loadQIdxForDataInValid & _T_93777; // @[AxiLoadQueue.scala 262:45:@39369.6]
  assign _T_93779 = _T_93778 | bypassRequest_14; // @[AxiLoadQueue.scala 262:78:@39370.6]
  assign _GEN_2092 = _T_93779 ? 1'h1 : dataKnown_14; // @[AxiLoadQueue.scala 262:99:@39371.6]
  assign _GEN_2093 = initBits_14 ? 1'h0 : _GEN_2092; // @[AxiLoadQueue.scala 260:25:@39364.4]
  assign _T_93783 = io_loadQIdxForDataIn == 32'hf; // @[AxiLoadQueue.scala 262:69:@39378.6]
  assign _T_93784 = io_loadQIdxForDataInValid & _T_93783; // @[AxiLoadQueue.scala 262:45:@39379.6]
  assign _T_93785 = _T_93784 | bypassRequest_15; // @[AxiLoadQueue.scala 262:78:@39380.6]
  assign _GEN_2094 = _T_93785 ? 1'h1 : dataKnown_15; // @[AxiLoadQueue.scala 262:99:@39381.6]
  assign _GEN_2095 = initBits_15 ? 1'h0 : _GEN_2094; // @[AxiLoadQueue.scala 260:25:@39374.4]
  assign _GEN_2096 = _T_93694 ? io_loadDataFromMem : dataQ_0; // @[AxiLoadQueue.scala 270:79:@39390.6]
  assign _GEN_2097 = bypassRequest_0 ? bypassVal_0 : _GEN_2096; // @[AxiLoadQueue.scala 268:32:@39384.4]
  assign _GEN_2098 = _T_93700 ? io_loadDataFromMem : dataQ_1; // @[AxiLoadQueue.scala 270:79:@39399.6]
  assign _GEN_2099 = bypassRequest_1 ? bypassVal_1 : _GEN_2098; // @[AxiLoadQueue.scala 268:32:@39393.4]
  assign _GEN_2100 = _T_93706 ? io_loadDataFromMem : dataQ_2; // @[AxiLoadQueue.scala 270:79:@39408.6]
  assign _GEN_2101 = bypassRequest_2 ? bypassVal_2 : _GEN_2100; // @[AxiLoadQueue.scala 268:32:@39402.4]
  assign _GEN_2102 = _T_93712 ? io_loadDataFromMem : dataQ_3; // @[AxiLoadQueue.scala 270:79:@39417.6]
  assign _GEN_2103 = bypassRequest_3 ? bypassVal_3 : _GEN_2102; // @[AxiLoadQueue.scala 268:32:@39411.4]
  assign _GEN_2104 = _T_93718 ? io_loadDataFromMem : dataQ_4; // @[AxiLoadQueue.scala 270:79:@39426.6]
  assign _GEN_2105 = bypassRequest_4 ? bypassVal_4 : _GEN_2104; // @[AxiLoadQueue.scala 268:32:@39420.4]
  assign _GEN_2106 = _T_93724 ? io_loadDataFromMem : dataQ_5; // @[AxiLoadQueue.scala 270:79:@39435.6]
  assign _GEN_2107 = bypassRequest_5 ? bypassVal_5 : _GEN_2106; // @[AxiLoadQueue.scala 268:32:@39429.4]
  assign _GEN_2108 = _T_93730 ? io_loadDataFromMem : dataQ_6; // @[AxiLoadQueue.scala 270:79:@39444.6]
  assign _GEN_2109 = bypassRequest_6 ? bypassVal_6 : _GEN_2108; // @[AxiLoadQueue.scala 268:32:@39438.4]
  assign _GEN_2110 = _T_93736 ? io_loadDataFromMem : dataQ_7; // @[AxiLoadQueue.scala 270:79:@39453.6]
  assign _GEN_2111 = bypassRequest_7 ? bypassVal_7 : _GEN_2110; // @[AxiLoadQueue.scala 268:32:@39447.4]
  assign _GEN_2112 = _T_93742 ? io_loadDataFromMem : dataQ_8; // @[AxiLoadQueue.scala 270:79:@39462.6]
  assign _GEN_2113 = bypassRequest_8 ? bypassVal_8 : _GEN_2112; // @[AxiLoadQueue.scala 268:32:@39456.4]
  assign _GEN_2114 = _T_93748 ? io_loadDataFromMem : dataQ_9; // @[AxiLoadQueue.scala 270:79:@39471.6]
  assign _GEN_2115 = bypassRequest_9 ? bypassVal_9 : _GEN_2114; // @[AxiLoadQueue.scala 268:32:@39465.4]
  assign _GEN_2116 = _T_93754 ? io_loadDataFromMem : dataQ_10; // @[AxiLoadQueue.scala 270:79:@39480.6]
  assign _GEN_2117 = bypassRequest_10 ? bypassVal_10 : _GEN_2116; // @[AxiLoadQueue.scala 268:32:@39474.4]
  assign _GEN_2118 = _T_93760 ? io_loadDataFromMem : dataQ_11; // @[AxiLoadQueue.scala 270:79:@39489.6]
  assign _GEN_2119 = bypassRequest_11 ? bypassVal_11 : _GEN_2118; // @[AxiLoadQueue.scala 268:32:@39483.4]
  assign _GEN_2120 = _T_93766 ? io_loadDataFromMem : dataQ_12; // @[AxiLoadQueue.scala 270:79:@39498.6]
  assign _GEN_2121 = bypassRequest_12 ? bypassVal_12 : _GEN_2120; // @[AxiLoadQueue.scala 268:32:@39492.4]
  assign _GEN_2122 = _T_93772 ? io_loadDataFromMem : dataQ_13; // @[AxiLoadQueue.scala 270:79:@39507.6]
  assign _GEN_2123 = bypassRequest_13 ? bypassVal_13 : _GEN_2122; // @[AxiLoadQueue.scala 268:32:@39501.4]
  assign _GEN_2124 = _T_93778 ? io_loadDataFromMem : dataQ_14; // @[AxiLoadQueue.scala 270:79:@39516.6]
  assign _GEN_2125 = bypassRequest_14 ? bypassVal_14 : _GEN_2124; // @[AxiLoadQueue.scala 268:32:@39510.4]
  assign _GEN_2126 = _T_93784 ? io_loadDataFromMem : dataQ_15; // @[AxiLoadQueue.scala 270:79:@39525.6]
  assign _GEN_2127 = bypassRequest_15 ? bypassVal_15 : _GEN_2126; // @[AxiLoadQueue.scala 268:32:@39519.4]
  assign entriesPorts_0_0 = portQ_0 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39529.4]
  assign entriesPorts_0_1 = portQ_1 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39531.4]
  assign entriesPorts_0_2 = portQ_2 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39533.4]
  assign entriesPorts_0_3 = portQ_3 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39535.4]
  assign entriesPorts_0_4 = portQ_4 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39537.4]
  assign entriesPorts_0_5 = portQ_5 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39539.4]
  assign entriesPorts_0_6 = portQ_6 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39541.4]
  assign entriesPorts_0_7 = portQ_7 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39543.4]
  assign entriesPorts_0_8 = portQ_8 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39545.4]
  assign entriesPorts_0_9 = portQ_9 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39547.4]
  assign entriesPorts_0_10 = portQ_10 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39549.4]
  assign entriesPorts_0_11 = portQ_11 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39551.4]
  assign entriesPorts_0_12 = portQ_12 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39553.4]
  assign entriesPorts_0_13 = portQ_13 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39555.4]
  assign entriesPorts_0_14 = portQ_14 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39557.4]
  assign entriesPorts_0_15 = portQ_15 == 1'h0; // @[AxiLoadQueue.scala 288:69:@39559.4]
  assign _T_94318 = addrKnown_0 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39563.4]
  assign _T_94319 = entriesPorts_0_0 & _T_94318; // @[AxiLoadQueue.scala 300:83:@39564.4]
  assign _T_94321 = addrKnown_1 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39565.4]
  assign _T_94322 = entriesPorts_0_1 & _T_94321; // @[AxiLoadQueue.scala 300:83:@39566.4]
  assign _T_94324 = addrKnown_2 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39567.4]
  assign _T_94325 = entriesPorts_0_2 & _T_94324; // @[AxiLoadQueue.scala 300:83:@39568.4]
  assign _T_94327 = addrKnown_3 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39569.4]
  assign _T_94328 = entriesPorts_0_3 & _T_94327; // @[AxiLoadQueue.scala 300:83:@39570.4]
  assign _T_94330 = addrKnown_4 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39571.4]
  assign _T_94331 = entriesPorts_0_4 & _T_94330; // @[AxiLoadQueue.scala 300:83:@39572.4]
  assign _T_94333 = addrKnown_5 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39573.4]
  assign _T_94334 = entriesPorts_0_5 & _T_94333; // @[AxiLoadQueue.scala 300:83:@39574.4]
  assign _T_94336 = addrKnown_6 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39575.4]
  assign _T_94337 = entriesPorts_0_6 & _T_94336; // @[AxiLoadQueue.scala 300:83:@39576.4]
  assign _T_94339 = addrKnown_7 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39577.4]
  assign _T_94340 = entriesPorts_0_7 & _T_94339; // @[AxiLoadQueue.scala 300:83:@39578.4]
  assign _T_94342 = addrKnown_8 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39579.4]
  assign _T_94343 = entriesPorts_0_8 & _T_94342; // @[AxiLoadQueue.scala 300:83:@39580.4]
  assign _T_94345 = addrKnown_9 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39581.4]
  assign _T_94346 = entriesPorts_0_9 & _T_94345; // @[AxiLoadQueue.scala 300:83:@39582.4]
  assign _T_94348 = addrKnown_10 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39583.4]
  assign _T_94349 = entriesPorts_0_10 & _T_94348; // @[AxiLoadQueue.scala 300:83:@39584.4]
  assign _T_94351 = addrKnown_11 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39585.4]
  assign _T_94352 = entriesPorts_0_11 & _T_94351; // @[AxiLoadQueue.scala 300:83:@39586.4]
  assign _T_94354 = addrKnown_12 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39587.4]
  assign _T_94355 = entriesPorts_0_12 & _T_94354; // @[AxiLoadQueue.scala 300:83:@39588.4]
  assign _T_94357 = addrKnown_13 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39589.4]
  assign _T_94358 = entriesPorts_0_13 & _T_94357; // @[AxiLoadQueue.scala 300:83:@39590.4]
  assign _T_94360 = addrKnown_14 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39591.4]
  assign _T_94361 = entriesPorts_0_14 & _T_94360; // @[AxiLoadQueue.scala 300:83:@39592.4]
  assign _T_94363 = addrKnown_15 == 1'h0; // @[AxiLoadQueue.scala 300:86:@39593.4]
  assign _T_94364 = entriesPorts_0_15 & _T_94363; // @[AxiLoadQueue.scala 300:83:@39594.4]
  assign _T_94447 = _T_94364 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39648.4]
  assign _T_94448 = _T_94361 ? 16'h4000 : _T_94447; // @[Mux.scala 31:69:@39649.4]
  assign _T_94449 = _T_94358 ? 16'h2000 : _T_94448; // @[Mux.scala 31:69:@39650.4]
  assign _T_94450 = _T_94355 ? 16'h1000 : _T_94449; // @[Mux.scala 31:69:@39651.4]
  assign _T_94451 = _T_94352 ? 16'h800 : _T_94450; // @[Mux.scala 31:69:@39652.4]
  assign _T_94452 = _T_94349 ? 16'h400 : _T_94451; // @[Mux.scala 31:69:@39653.4]
  assign _T_94453 = _T_94346 ? 16'h200 : _T_94452; // @[Mux.scala 31:69:@39654.4]
  assign _T_94454 = _T_94343 ? 16'h100 : _T_94453; // @[Mux.scala 31:69:@39655.4]
  assign _T_94455 = _T_94340 ? 16'h80 : _T_94454; // @[Mux.scala 31:69:@39656.4]
  assign _T_94456 = _T_94337 ? 16'h40 : _T_94455; // @[Mux.scala 31:69:@39657.4]
  assign _T_94457 = _T_94334 ? 16'h20 : _T_94456; // @[Mux.scala 31:69:@39658.4]
  assign _T_94458 = _T_94331 ? 16'h10 : _T_94457; // @[Mux.scala 31:69:@39659.4]
  assign _T_94459 = _T_94328 ? 16'h8 : _T_94458; // @[Mux.scala 31:69:@39660.4]
  assign _T_94460 = _T_94325 ? 16'h4 : _T_94459; // @[Mux.scala 31:69:@39661.4]
  assign _T_94461 = _T_94322 ? 16'h2 : _T_94460; // @[Mux.scala 31:69:@39662.4]
  assign _T_94462 = _T_94319 ? 16'h1 : _T_94461; // @[Mux.scala 31:69:@39663.4]
  assign _T_94463 = _T_94462[0]; // @[OneHot.scala 66:30:@39664.4]
  assign _T_94464 = _T_94462[1]; // @[OneHot.scala 66:30:@39665.4]
  assign _T_94465 = _T_94462[2]; // @[OneHot.scala 66:30:@39666.4]
  assign _T_94466 = _T_94462[3]; // @[OneHot.scala 66:30:@39667.4]
  assign _T_94467 = _T_94462[4]; // @[OneHot.scala 66:30:@39668.4]
  assign _T_94468 = _T_94462[5]; // @[OneHot.scala 66:30:@39669.4]
  assign _T_94469 = _T_94462[6]; // @[OneHot.scala 66:30:@39670.4]
  assign _T_94470 = _T_94462[7]; // @[OneHot.scala 66:30:@39671.4]
  assign _T_94471 = _T_94462[8]; // @[OneHot.scala 66:30:@39672.4]
  assign _T_94472 = _T_94462[9]; // @[OneHot.scala 66:30:@39673.4]
  assign _T_94473 = _T_94462[10]; // @[OneHot.scala 66:30:@39674.4]
  assign _T_94474 = _T_94462[11]; // @[OneHot.scala 66:30:@39675.4]
  assign _T_94475 = _T_94462[12]; // @[OneHot.scala 66:30:@39676.4]
  assign _T_94476 = _T_94462[13]; // @[OneHot.scala 66:30:@39677.4]
  assign _T_94477 = _T_94462[14]; // @[OneHot.scala 66:30:@39678.4]
  assign _T_94478 = _T_94462[15]; // @[OneHot.scala 66:30:@39679.4]
  assign _T_94519 = _T_94319 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39697.4]
  assign _T_94520 = _T_94364 ? 16'h4000 : _T_94519; // @[Mux.scala 31:69:@39698.4]
  assign _T_94521 = _T_94361 ? 16'h2000 : _T_94520; // @[Mux.scala 31:69:@39699.4]
  assign _T_94522 = _T_94358 ? 16'h1000 : _T_94521; // @[Mux.scala 31:69:@39700.4]
  assign _T_94523 = _T_94355 ? 16'h800 : _T_94522; // @[Mux.scala 31:69:@39701.4]
  assign _T_94524 = _T_94352 ? 16'h400 : _T_94523; // @[Mux.scala 31:69:@39702.4]
  assign _T_94525 = _T_94349 ? 16'h200 : _T_94524; // @[Mux.scala 31:69:@39703.4]
  assign _T_94526 = _T_94346 ? 16'h100 : _T_94525; // @[Mux.scala 31:69:@39704.4]
  assign _T_94527 = _T_94343 ? 16'h80 : _T_94526; // @[Mux.scala 31:69:@39705.4]
  assign _T_94528 = _T_94340 ? 16'h40 : _T_94527; // @[Mux.scala 31:69:@39706.4]
  assign _T_94529 = _T_94337 ? 16'h20 : _T_94528; // @[Mux.scala 31:69:@39707.4]
  assign _T_94530 = _T_94334 ? 16'h10 : _T_94529; // @[Mux.scala 31:69:@39708.4]
  assign _T_94531 = _T_94331 ? 16'h8 : _T_94530; // @[Mux.scala 31:69:@39709.4]
  assign _T_94532 = _T_94328 ? 16'h4 : _T_94531; // @[Mux.scala 31:69:@39710.4]
  assign _T_94533 = _T_94325 ? 16'h2 : _T_94532; // @[Mux.scala 31:69:@39711.4]
  assign _T_94534 = _T_94322 ? 16'h1 : _T_94533; // @[Mux.scala 31:69:@39712.4]
  assign _T_94535 = _T_94534[0]; // @[OneHot.scala 66:30:@39713.4]
  assign _T_94536 = _T_94534[1]; // @[OneHot.scala 66:30:@39714.4]
  assign _T_94537 = _T_94534[2]; // @[OneHot.scala 66:30:@39715.4]
  assign _T_94538 = _T_94534[3]; // @[OneHot.scala 66:30:@39716.4]
  assign _T_94539 = _T_94534[4]; // @[OneHot.scala 66:30:@39717.4]
  assign _T_94540 = _T_94534[5]; // @[OneHot.scala 66:30:@39718.4]
  assign _T_94541 = _T_94534[6]; // @[OneHot.scala 66:30:@39719.4]
  assign _T_94542 = _T_94534[7]; // @[OneHot.scala 66:30:@39720.4]
  assign _T_94543 = _T_94534[8]; // @[OneHot.scala 66:30:@39721.4]
  assign _T_94544 = _T_94534[9]; // @[OneHot.scala 66:30:@39722.4]
  assign _T_94545 = _T_94534[10]; // @[OneHot.scala 66:30:@39723.4]
  assign _T_94546 = _T_94534[11]; // @[OneHot.scala 66:30:@39724.4]
  assign _T_94547 = _T_94534[12]; // @[OneHot.scala 66:30:@39725.4]
  assign _T_94548 = _T_94534[13]; // @[OneHot.scala 66:30:@39726.4]
  assign _T_94549 = _T_94534[14]; // @[OneHot.scala 66:30:@39727.4]
  assign _T_94550 = _T_94534[15]; // @[OneHot.scala 66:30:@39728.4]
  assign _T_94591 = _T_94322 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39746.4]
  assign _T_94592 = _T_94319 ? 16'h4000 : _T_94591; // @[Mux.scala 31:69:@39747.4]
  assign _T_94593 = _T_94364 ? 16'h2000 : _T_94592; // @[Mux.scala 31:69:@39748.4]
  assign _T_94594 = _T_94361 ? 16'h1000 : _T_94593; // @[Mux.scala 31:69:@39749.4]
  assign _T_94595 = _T_94358 ? 16'h800 : _T_94594; // @[Mux.scala 31:69:@39750.4]
  assign _T_94596 = _T_94355 ? 16'h400 : _T_94595; // @[Mux.scala 31:69:@39751.4]
  assign _T_94597 = _T_94352 ? 16'h200 : _T_94596; // @[Mux.scala 31:69:@39752.4]
  assign _T_94598 = _T_94349 ? 16'h100 : _T_94597; // @[Mux.scala 31:69:@39753.4]
  assign _T_94599 = _T_94346 ? 16'h80 : _T_94598; // @[Mux.scala 31:69:@39754.4]
  assign _T_94600 = _T_94343 ? 16'h40 : _T_94599; // @[Mux.scala 31:69:@39755.4]
  assign _T_94601 = _T_94340 ? 16'h20 : _T_94600; // @[Mux.scala 31:69:@39756.4]
  assign _T_94602 = _T_94337 ? 16'h10 : _T_94601; // @[Mux.scala 31:69:@39757.4]
  assign _T_94603 = _T_94334 ? 16'h8 : _T_94602; // @[Mux.scala 31:69:@39758.4]
  assign _T_94604 = _T_94331 ? 16'h4 : _T_94603; // @[Mux.scala 31:69:@39759.4]
  assign _T_94605 = _T_94328 ? 16'h2 : _T_94604; // @[Mux.scala 31:69:@39760.4]
  assign _T_94606 = _T_94325 ? 16'h1 : _T_94605; // @[Mux.scala 31:69:@39761.4]
  assign _T_94607 = _T_94606[0]; // @[OneHot.scala 66:30:@39762.4]
  assign _T_94608 = _T_94606[1]; // @[OneHot.scala 66:30:@39763.4]
  assign _T_94609 = _T_94606[2]; // @[OneHot.scala 66:30:@39764.4]
  assign _T_94610 = _T_94606[3]; // @[OneHot.scala 66:30:@39765.4]
  assign _T_94611 = _T_94606[4]; // @[OneHot.scala 66:30:@39766.4]
  assign _T_94612 = _T_94606[5]; // @[OneHot.scala 66:30:@39767.4]
  assign _T_94613 = _T_94606[6]; // @[OneHot.scala 66:30:@39768.4]
  assign _T_94614 = _T_94606[7]; // @[OneHot.scala 66:30:@39769.4]
  assign _T_94615 = _T_94606[8]; // @[OneHot.scala 66:30:@39770.4]
  assign _T_94616 = _T_94606[9]; // @[OneHot.scala 66:30:@39771.4]
  assign _T_94617 = _T_94606[10]; // @[OneHot.scala 66:30:@39772.4]
  assign _T_94618 = _T_94606[11]; // @[OneHot.scala 66:30:@39773.4]
  assign _T_94619 = _T_94606[12]; // @[OneHot.scala 66:30:@39774.4]
  assign _T_94620 = _T_94606[13]; // @[OneHot.scala 66:30:@39775.4]
  assign _T_94621 = _T_94606[14]; // @[OneHot.scala 66:30:@39776.4]
  assign _T_94622 = _T_94606[15]; // @[OneHot.scala 66:30:@39777.4]
  assign _T_94663 = _T_94325 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39795.4]
  assign _T_94664 = _T_94322 ? 16'h4000 : _T_94663; // @[Mux.scala 31:69:@39796.4]
  assign _T_94665 = _T_94319 ? 16'h2000 : _T_94664; // @[Mux.scala 31:69:@39797.4]
  assign _T_94666 = _T_94364 ? 16'h1000 : _T_94665; // @[Mux.scala 31:69:@39798.4]
  assign _T_94667 = _T_94361 ? 16'h800 : _T_94666; // @[Mux.scala 31:69:@39799.4]
  assign _T_94668 = _T_94358 ? 16'h400 : _T_94667; // @[Mux.scala 31:69:@39800.4]
  assign _T_94669 = _T_94355 ? 16'h200 : _T_94668; // @[Mux.scala 31:69:@39801.4]
  assign _T_94670 = _T_94352 ? 16'h100 : _T_94669; // @[Mux.scala 31:69:@39802.4]
  assign _T_94671 = _T_94349 ? 16'h80 : _T_94670; // @[Mux.scala 31:69:@39803.4]
  assign _T_94672 = _T_94346 ? 16'h40 : _T_94671; // @[Mux.scala 31:69:@39804.4]
  assign _T_94673 = _T_94343 ? 16'h20 : _T_94672; // @[Mux.scala 31:69:@39805.4]
  assign _T_94674 = _T_94340 ? 16'h10 : _T_94673; // @[Mux.scala 31:69:@39806.4]
  assign _T_94675 = _T_94337 ? 16'h8 : _T_94674; // @[Mux.scala 31:69:@39807.4]
  assign _T_94676 = _T_94334 ? 16'h4 : _T_94675; // @[Mux.scala 31:69:@39808.4]
  assign _T_94677 = _T_94331 ? 16'h2 : _T_94676; // @[Mux.scala 31:69:@39809.4]
  assign _T_94678 = _T_94328 ? 16'h1 : _T_94677; // @[Mux.scala 31:69:@39810.4]
  assign _T_94679 = _T_94678[0]; // @[OneHot.scala 66:30:@39811.4]
  assign _T_94680 = _T_94678[1]; // @[OneHot.scala 66:30:@39812.4]
  assign _T_94681 = _T_94678[2]; // @[OneHot.scala 66:30:@39813.4]
  assign _T_94682 = _T_94678[3]; // @[OneHot.scala 66:30:@39814.4]
  assign _T_94683 = _T_94678[4]; // @[OneHot.scala 66:30:@39815.4]
  assign _T_94684 = _T_94678[5]; // @[OneHot.scala 66:30:@39816.4]
  assign _T_94685 = _T_94678[6]; // @[OneHot.scala 66:30:@39817.4]
  assign _T_94686 = _T_94678[7]; // @[OneHot.scala 66:30:@39818.4]
  assign _T_94687 = _T_94678[8]; // @[OneHot.scala 66:30:@39819.4]
  assign _T_94688 = _T_94678[9]; // @[OneHot.scala 66:30:@39820.4]
  assign _T_94689 = _T_94678[10]; // @[OneHot.scala 66:30:@39821.4]
  assign _T_94690 = _T_94678[11]; // @[OneHot.scala 66:30:@39822.4]
  assign _T_94691 = _T_94678[12]; // @[OneHot.scala 66:30:@39823.4]
  assign _T_94692 = _T_94678[13]; // @[OneHot.scala 66:30:@39824.4]
  assign _T_94693 = _T_94678[14]; // @[OneHot.scala 66:30:@39825.4]
  assign _T_94694 = _T_94678[15]; // @[OneHot.scala 66:30:@39826.4]
  assign _T_94735 = _T_94328 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39844.4]
  assign _T_94736 = _T_94325 ? 16'h4000 : _T_94735; // @[Mux.scala 31:69:@39845.4]
  assign _T_94737 = _T_94322 ? 16'h2000 : _T_94736; // @[Mux.scala 31:69:@39846.4]
  assign _T_94738 = _T_94319 ? 16'h1000 : _T_94737; // @[Mux.scala 31:69:@39847.4]
  assign _T_94739 = _T_94364 ? 16'h800 : _T_94738; // @[Mux.scala 31:69:@39848.4]
  assign _T_94740 = _T_94361 ? 16'h400 : _T_94739; // @[Mux.scala 31:69:@39849.4]
  assign _T_94741 = _T_94358 ? 16'h200 : _T_94740; // @[Mux.scala 31:69:@39850.4]
  assign _T_94742 = _T_94355 ? 16'h100 : _T_94741; // @[Mux.scala 31:69:@39851.4]
  assign _T_94743 = _T_94352 ? 16'h80 : _T_94742; // @[Mux.scala 31:69:@39852.4]
  assign _T_94744 = _T_94349 ? 16'h40 : _T_94743; // @[Mux.scala 31:69:@39853.4]
  assign _T_94745 = _T_94346 ? 16'h20 : _T_94744; // @[Mux.scala 31:69:@39854.4]
  assign _T_94746 = _T_94343 ? 16'h10 : _T_94745; // @[Mux.scala 31:69:@39855.4]
  assign _T_94747 = _T_94340 ? 16'h8 : _T_94746; // @[Mux.scala 31:69:@39856.4]
  assign _T_94748 = _T_94337 ? 16'h4 : _T_94747; // @[Mux.scala 31:69:@39857.4]
  assign _T_94749 = _T_94334 ? 16'h2 : _T_94748; // @[Mux.scala 31:69:@39858.4]
  assign _T_94750 = _T_94331 ? 16'h1 : _T_94749; // @[Mux.scala 31:69:@39859.4]
  assign _T_94751 = _T_94750[0]; // @[OneHot.scala 66:30:@39860.4]
  assign _T_94752 = _T_94750[1]; // @[OneHot.scala 66:30:@39861.4]
  assign _T_94753 = _T_94750[2]; // @[OneHot.scala 66:30:@39862.4]
  assign _T_94754 = _T_94750[3]; // @[OneHot.scala 66:30:@39863.4]
  assign _T_94755 = _T_94750[4]; // @[OneHot.scala 66:30:@39864.4]
  assign _T_94756 = _T_94750[5]; // @[OneHot.scala 66:30:@39865.4]
  assign _T_94757 = _T_94750[6]; // @[OneHot.scala 66:30:@39866.4]
  assign _T_94758 = _T_94750[7]; // @[OneHot.scala 66:30:@39867.4]
  assign _T_94759 = _T_94750[8]; // @[OneHot.scala 66:30:@39868.4]
  assign _T_94760 = _T_94750[9]; // @[OneHot.scala 66:30:@39869.4]
  assign _T_94761 = _T_94750[10]; // @[OneHot.scala 66:30:@39870.4]
  assign _T_94762 = _T_94750[11]; // @[OneHot.scala 66:30:@39871.4]
  assign _T_94763 = _T_94750[12]; // @[OneHot.scala 66:30:@39872.4]
  assign _T_94764 = _T_94750[13]; // @[OneHot.scala 66:30:@39873.4]
  assign _T_94765 = _T_94750[14]; // @[OneHot.scala 66:30:@39874.4]
  assign _T_94766 = _T_94750[15]; // @[OneHot.scala 66:30:@39875.4]
  assign _T_94807 = _T_94331 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39893.4]
  assign _T_94808 = _T_94328 ? 16'h4000 : _T_94807; // @[Mux.scala 31:69:@39894.4]
  assign _T_94809 = _T_94325 ? 16'h2000 : _T_94808; // @[Mux.scala 31:69:@39895.4]
  assign _T_94810 = _T_94322 ? 16'h1000 : _T_94809; // @[Mux.scala 31:69:@39896.4]
  assign _T_94811 = _T_94319 ? 16'h800 : _T_94810; // @[Mux.scala 31:69:@39897.4]
  assign _T_94812 = _T_94364 ? 16'h400 : _T_94811; // @[Mux.scala 31:69:@39898.4]
  assign _T_94813 = _T_94361 ? 16'h200 : _T_94812; // @[Mux.scala 31:69:@39899.4]
  assign _T_94814 = _T_94358 ? 16'h100 : _T_94813; // @[Mux.scala 31:69:@39900.4]
  assign _T_94815 = _T_94355 ? 16'h80 : _T_94814; // @[Mux.scala 31:69:@39901.4]
  assign _T_94816 = _T_94352 ? 16'h40 : _T_94815; // @[Mux.scala 31:69:@39902.4]
  assign _T_94817 = _T_94349 ? 16'h20 : _T_94816; // @[Mux.scala 31:69:@39903.4]
  assign _T_94818 = _T_94346 ? 16'h10 : _T_94817; // @[Mux.scala 31:69:@39904.4]
  assign _T_94819 = _T_94343 ? 16'h8 : _T_94818; // @[Mux.scala 31:69:@39905.4]
  assign _T_94820 = _T_94340 ? 16'h4 : _T_94819; // @[Mux.scala 31:69:@39906.4]
  assign _T_94821 = _T_94337 ? 16'h2 : _T_94820; // @[Mux.scala 31:69:@39907.4]
  assign _T_94822 = _T_94334 ? 16'h1 : _T_94821; // @[Mux.scala 31:69:@39908.4]
  assign _T_94823 = _T_94822[0]; // @[OneHot.scala 66:30:@39909.4]
  assign _T_94824 = _T_94822[1]; // @[OneHot.scala 66:30:@39910.4]
  assign _T_94825 = _T_94822[2]; // @[OneHot.scala 66:30:@39911.4]
  assign _T_94826 = _T_94822[3]; // @[OneHot.scala 66:30:@39912.4]
  assign _T_94827 = _T_94822[4]; // @[OneHot.scala 66:30:@39913.4]
  assign _T_94828 = _T_94822[5]; // @[OneHot.scala 66:30:@39914.4]
  assign _T_94829 = _T_94822[6]; // @[OneHot.scala 66:30:@39915.4]
  assign _T_94830 = _T_94822[7]; // @[OneHot.scala 66:30:@39916.4]
  assign _T_94831 = _T_94822[8]; // @[OneHot.scala 66:30:@39917.4]
  assign _T_94832 = _T_94822[9]; // @[OneHot.scala 66:30:@39918.4]
  assign _T_94833 = _T_94822[10]; // @[OneHot.scala 66:30:@39919.4]
  assign _T_94834 = _T_94822[11]; // @[OneHot.scala 66:30:@39920.4]
  assign _T_94835 = _T_94822[12]; // @[OneHot.scala 66:30:@39921.4]
  assign _T_94836 = _T_94822[13]; // @[OneHot.scala 66:30:@39922.4]
  assign _T_94837 = _T_94822[14]; // @[OneHot.scala 66:30:@39923.4]
  assign _T_94838 = _T_94822[15]; // @[OneHot.scala 66:30:@39924.4]
  assign _T_94879 = _T_94334 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39942.4]
  assign _T_94880 = _T_94331 ? 16'h4000 : _T_94879; // @[Mux.scala 31:69:@39943.4]
  assign _T_94881 = _T_94328 ? 16'h2000 : _T_94880; // @[Mux.scala 31:69:@39944.4]
  assign _T_94882 = _T_94325 ? 16'h1000 : _T_94881; // @[Mux.scala 31:69:@39945.4]
  assign _T_94883 = _T_94322 ? 16'h800 : _T_94882; // @[Mux.scala 31:69:@39946.4]
  assign _T_94884 = _T_94319 ? 16'h400 : _T_94883; // @[Mux.scala 31:69:@39947.4]
  assign _T_94885 = _T_94364 ? 16'h200 : _T_94884; // @[Mux.scala 31:69:@39948.4]
  assign _T_94886 = _T_94361 ? 16'h100 : _T_94885; // @[Mux.scala 31:69:@39949.4]
  assign _T_94887 = _T_94358 ? 16'h80 : _T_94886; // @[Mux.scala 31:69:@39950.4]
  assign _T_94888 = _T_94355 ? 16'h40 : _T_94887; // @[Mux.scala 31:69:@39951.4]
  assign _T_94889 = _T_94352 ? 16'h20 : _T_94888; // @[Mux.scala 31:69:@39952.4]
  assign _T_94890 = _T_94349 ? 16'h10 : _T_94889; // @[Mux.scala 31:69:@39953.4]
  assign _T_94891 = _T_94346 ? 16'h8 : _T_94890; // @[Mux.scala 31:69:@39954.4]
  assign _T_94892 = _T_94343 ? 16'h4 : _T_94891; // @[Mux.scala 31:69:@39955.4]
  assign _T_94893 = _T_94340 ? 16'h2 : _T_94892; // @[Mux.scala 31:69:@39956.4]
  assign _T_94894 = _T_94337 ? 16'h1 : _T_94893; // @[Mux.scala 31:69:@39957.4]
  assign _T_94895 = _T_94894[0]; // @[OneHot.scala 66:30:@39958.4]
  assign _T_94896 = _T_94894[1]; // @[OneHot.scala 66:30:@39959.4]
  assign _T_94897 = _T_94894[2]; // @[OneHot.scala 66:30:@39960.4]
  assign _T_94898 = _T_94894[3]; // @[OneHot.scala 66:30:@39961.4]
  assign _T_94899 = _T_94894[4]; // @[OneHot.scala 66:30:@39962.4]
  assign _T_94900 = _T_94894[5]; // @[OneHot.scala 66:30:@39963.4]
  assign _T_94901 = _T_94894[6]; // @[OneHot.scala 66:30:@39964.4]
  assign _T_94902 = _T_94894[7]; // @[OneHot.scala 66:30:@39965.4]
  assign _T_94903 = _T_94894[8]; // @[OneHot.scala 66:30:@39966.4]
  assign _T_94904 = _T_94894[9]; // @[OneHot.scala 66:30:@39967.4]
  assign _T_94905 = _T_94894[10]; // @[OneHot.scala 66:30:@39968.4]
  assign _T_94906 = _T_94894[11]; // @[OneHot.scala 66:30:@39969.4]
  assign _T_94907 = _T_94894[12]; // @[OneHot.scala 66:30:@39970.4]
  assign _T_94908 = _T_94894[13]; // @[OneHot.scala 66:30:@39971.4]
  assign _T_94909 = _T_94894[14]; // @[OneHot.scala 66:30:@39972.4]
  assign _T_94910 = _T_94894[15]; // @[OneHot.scala 66:30:@39973.4]
  assign _T_94951 = _T_94337 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@39991.4]
  assign _T_94952 = _T_94334 ? 16'h4000 : _T_94951; // @[Mux.scala 31:69:@39992.4]
  assign _T_94953 = _T_94331 ? 16'h2000 : _T_94952; // @[Mux.scala 31:69:@39993.4]
  assign _T_94954 = _T_94328 ? 16'h1000 : _T_94953; // @[Mux.scala 31:69:@39994.4]
  assign _T_94955 = _T_94325 ? 16'h800 : _T_94954; // @[Mux.scala 31:69:@39995.4]
  assign _T_94956 = _T_94322 ? 16'h400 : _T_94955; // @[Mux.scala 31:69:@39996.4]
  assign _T_94957 = _T_94319 ? 16'h200 : _T_94956; // @[Mux.scala 31:69:@39997.4]
  assign _T_94958 = _T_94364 ? 16'h100 : _T_94957; // @[Mux.scala 31:69:@39998.4]
  assign _T_94959 = _T_94361 ? 16'h80 : _T_94958; // @[Mux.scala 31:69:@39999.4]
  assign _T_94960 = _T_94358 ? 16'h40 : _T_94959; // @[Mux.scala 31:69:@40000.4]
  assign _T_94961 = _T_94355 ? 16'h20 : _T_94960; // @[Mux.scala 31:69:@40001.4]
  assign _T_94962 = _T_94352 ? 16'h10 : _T_94961; // @[Mux.scala 31:69:@40002.4]
  assign _T_94963 = _T_94349 ? 16'h8 : _T_94962; // @[Mux.scala 31:69:@40003.4]
  assign _T_94964 = _T_94346 ? 16'h4 : _T_94963; // @[Mux.scala 31:69:@40004.4]
  assign _T_94965 = _T_94343 ? 16'h2 : _T_94964; // @[Mux.scala 31:69:@40005.4]
  assign _T_94966 = _T_94340 ? 16'h1 : _T_94965; // @[Mux.scala 31:69:@40006.4]
  assign _T_94967 = _T_94966[0]; // @[OneHot.scala 66:30:@40007.4]
  assign _T_94968 = _T_94966[1]; // @[OneHot.scala 66:30:@40008.4]
  assign _T_94969 = _T_94966[2]; // @[OneHot.scala 66:30:@40009.4]
  assign _T_94970 = _T_94966[3]; // @[OneHot.scala 66:30:@40010.4]
  assign _T_94971 = _T_94966[4]; // @[OneHot.scala 66:30:@40011.4]
  assign _T_94972 = _T_94966[5]; // @[OneHot.scala 66:30:@40012.4]
  assign _T_94973 = _T_94966[6]; // @[OneHot.scala 66:30:@40013.4]
  assign _T_94974 = _T_94966[7]; // @[OneHot.scala 66:30:@40014.4]
  assign _T_94975 = _T_94966[8]; // @[OneHot.scala 66:30:@40015.4]
  assign _T_94976 = _T_94966[9]; // @[OneHot.scala 66:30:@40016.4]
  assign _T_94977 = _T_94966[10]; // @[OneHot.scala 66:30:@40017.4]
  assign _T_94978 = _T_94966[11]; // @[OneHot.scala 66:30:@40018.4]
  assign _T_94979 = _T_94966[12]; // @[OneHot.scala 66:30:@40019.4]
  assign _T_94980 = _T_94966[13]; // @[OneHot.scala 66:30:@40020.4]
  assign _T_94981 = _T_94966[14]; // @[OneHot.scala 66:30:@40021.4]
  assign _T_94982 = _T_94966[15]; // @[OneHot.scala 66:30:@40022.4]
  assign _T_95023 = _T_94340 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40040.4]
  assign _T_95024 = _T_94337 ? 16'h4000 : _T_95023; // @[Mux.scala 31:69:@40041.4]
  assign _T_95025 = _T_94334 ? 16'h2000 : _T_95024; // @[Mux.scala 31:69:@40042.4]
  assign _T_95026 = _T_94331 ? 16'h1000 : _T_95025; // @[Mux.scala 31:69:@40043.4]
  assign _T_95027 = _T_94328 ? 16'h800 : _T_95026; // @[Mux.scala 31:69:@40044.4]
  assign _T_95028 = _T_94325 ? 16'h400 : _T_95027; // @[Mux.scala 31:69:@40045.4]
  assign _T_95029 = _T_94322 ? 16'h200 : _T_95028; // @[Mux.scala 31:69:@40046.4]
  assign _T_95030 = _T_94319 ? 16'h100 : _T_95029; // @[Mux.scala 31:69:@40047.4]
  assign _T_95031 = _T_94364 ? 16'h80 : _T_95030; // @[Mux.scala 31:69:@40048.4]
  assign _T_95032 = _T_94361 ? 16'h40 : _T_95031; // @[Mux.scala 31:69:@40049.4]
  assign _T_95033 = _T_94358 ? 16'h20 : _T_95032; // @[Mux.scala 31:69:@40050.4]
  assign _T_95034 = _T_94355 ? 16'h10 : _T_95033; // @[Mux.scala 31:69:@40051.4]
  assign _T_95035 = _T_94352 ? 16'h8 : _T_95034; // @[Mux.scala 31:69:@40052.4]
  assign _T_95036 = _T_94349 ? 16'h4 : _T_95035; // @[Mux.scala 31:69:@40053.4]
  assign _T_95037 = _T_94346 ? 16'h2 : _T_95036; // @[Mux.scala 31:69:@40054.4]
  assign _T_95038 = _T_94343 ? 16'h1 : _T_95037; // @[Mux.scala 31:69:@40055.4]
  assign _T_95039 = _T_95038[0]; // @[OneHot.scala 66:30:@40056.4]
  assign _T_95040 = _T_95038[1]; // @[OneHot.scala 66:30:@40057.4]
  assign _T_95041 = _T_95038[2]; // @[OneHot.scala 66:30:@40058.4]
  assign _T_95042 = _T_95038[3]; // @[OneHot.scala 66:30:@40059.4]
  assign _T_95043 = _T_95038[4]; // @[OneHot.scala 66:30:@40060.4]
  assign _T_95044 = _T_95038[5]; // @[OneHot.scala 66:30:@40061.4]
  assign _T_95045 = _T_95038[6]; // @[OneHot.scala 66:30:@40062.4]
  assign _T_95046 = _T_95038[7]; // @[OneHot.scala 66:30:@40063.4]
  assign _T_95047 = _T_95038[8]; // @[OneHot.scala 66:30:@40064.4]
  assign _T_95048 = _T_95038[9]; // @[OneHot.scala 66:30:@40065.4]
  assign _T_95049 = _T_95038[10]; // @[OneHot.scala 66:30:@40066.4]
  assign _T_95050 = _T_95038[11]; // @[OneHot.scala 66:30:@40067.4]
  assign _T_95051 = _T_95038[12]; // @[OneHot.scala 66:30:@40068.4]
  assign _T_95052 = _T_95038[13]; // @[OneHot.scala 66:30:@40069.4]
  assign _T_95053 = _T_95038[14]; // @[OneHot.scala 66:30:@40070.4]
  assign _T_95054 = _T_95038[15]; // @[OneHot.scala 66:30:@40071.4]
  assign _T_95095 = _T_94343 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40089.4]
  assign _T_95096 = _T_94340 ? 16'h4000 : _T_95095; // @[Mux.scala 31:69:@40090.4]
  assign _T_95097 = _T_94337 ? 16'h2000 : _T_95096; // @[Mux.scala 31:69:@40091.4]
  assign _T_95098 = _T_94334 ? 16'h1000 : _T_95097; // @[Mux.scala 31:69:@40092.4]
  assign _T_95099 = _T_94331 ? 16'h800 : _T_95098; // @[Mux.scala 31:69:@40093.4]
  assign _T_95100 = _T_94328 ? 16'h400 : _T_95099; // @[Mux.scala 31:69:@40094.4]
  assign _T_95101 = _T_94325 ? 16'h200 : _T_95100; // @[Mux.scala 31:69:@40095.4]
  assign _T_95102 = _T_94322 ? 16'h100 : _T_95101; // @[Mux.scala 31:69:@40096.4]
  assign _T_95103 = _T_94319 ? 16'h80 : _T_95102; // @[Mux.scala 31:69:@40097.4]
  assign _T_95104 = _T_94364 ? 16'h40 : _T_95103; // @[Mux.scala 31:69:@40098.4]
  assign _T_95105 = _T_94361 ? 16'h20 : _T_95104; // @[Mux.scala 31:69:@40099.4]
  assign _T_95106 = _T_94358 ? 16'h10 : _T_95105; // @[Mux.scala 31:69:@40100.4]
  assign _T_95107 = _T_94355 ? 16'h8 : _T_95106; // @[Mux.scala 31:69:@40101.4]
  assign _T_95108 = _T_94352 ? 16'h4 : _T_95107; // @[Mux.scala 31:69:@40102.4]
  assign _T_95109 = _T_94349 ? 16'h2 : _T_95108; // @[Mux.scala 31:69:@40103.4]
  assign _T_95110 = _T_94346 ? 16'h1 : _T_95109; // @[Mux.scala 31:69:@40104.4]
  assign _T_95111 = _T_95110[0]; // @[OneHot.scala 66:30:@40105.4]
  assign _T_95112 = _T_95110[1]; // @[OneHot.scala 66:30:@40106.4]
  assign _T_95113 = _T_95110[2]; // @[OneHot.scala 66:30:@40107.4]
  assign _T_95114 = _T_95110[3]; // @[OneHot.scala 66:30:@40108.4]
  assign _T_95115 = _T_95110[4]; // @[OneHot.scala 66:30:@40109.4]
  assign _T_95116 = _T_95110[5]; // @[OneHot.scala 66:30:@40110.4]
  assign _T_95117 = _T_95110[6]; // @[OneHot.scala 66:30:@40111.4]
  assign _T_95118 = _T_95110[7]; // @[OneHot.scala 66:30:@40112.4]
  assign _T_95119 = _T_95110[8]; // @[OneHot.scala 66:30:@40113.4]
  assign _T_95120 = _T_95110[9]; // @[OneHot.scala 66:30:@40114.4]
  assign _T_95121 = _T_95110[10]; // @[OneHot.scala 66:30:@40115.4]
  assign _T_95122 = _T_95110[11]; // @[OneHot.scala 66:30:@40116.4]
  assign _T_95123 = _T_95110[12]; // @[OneHot.scala 66:30:@40117.4]
  assign _T_95124 = _T_95110[13]; // @[OneHot.scala 66:30:@40118.4]
  assign _T_95125 = _T_95110[14]; // @[OneHot.scala 66:30:@40119.4]
  assign _T_95126 = _T_95110[15]; // @[OneHot.scala 66:30:@40120.4]
  assign _T_95167 = _T_94346 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40138.4]
  assign _T_95168 = _T_94343 ? 16'h4000 : _T_95167; // @[Mux.scala 31:69:@40139.4]
  assign _T_95169 = _T_94340 ? 16'h2000 : _T_95168; // @[Mux.scala 31:69:@40140.4]
  assign _T_95170 = _T_94337 ? 16'h1000 : _T_95169; // @[Mux.scala 31:69:@40141.4]
  assign _T_95171 = _T_94334 ? 16'h800 : _T_95170; // @[Mux.scala 31:69:@40142.4]
  assign _T_95172 = _T_94331 ? 16'h400 : _T_95171; // @[Mux.scala 31:69:@40143.4]
  assign _T_95173 = _T_94328 ? 16'h200 : _T_95172; // @[Mux.scala 31:69:@40144.4]
  assign _T_95174 = _T_94325 ? 16'h100 : _T_95173; // @[Mux.scala 31:69:@40145.4]
  assign _T_95175 = _T_94322 ? 16'h80 : _T_95174; // @[Mux.scala 31:69:@40146.4]
  assign _T_95176 = _T_94319 ? 16'h40 : _T_95175; // @[Mux.scala 31:69:@40147.4]
  assign _T_95177 = _T_94364 ? 16'h20 : _T_95176; // @[Mux.scala 31:69:@40148.4]
  assign _T_95178 = _T_94361 ? 16'h10 : _T_95177; // @[Mux.scala 31:69:@40149.4]
  assign _T_95179 = _T_94358 ? 16'h8 : _T_95178; // @[Mux.scala 31:69:@40150.4]
  assign _T_95180 = _T_94355 ? 16'h4 : _T_95179; // @[Mux.scala 31:69:@40151.4]
  assign _T_95181 = _T_94352 ? 16'h2 : _T_95180; // @[Mux.scala 31:69:@40152.4]
  assign _T_95182 = _T_94349 ? 16'h1 : _T_95181; // @[Mux.scala 31:69:@40153.4]
  assign _T_95183 = _T_95182[0]; // @[OneHot.scala 66:30:@40154.4]
  assign _T_95184 = _T_95182[1]; // @[OneHot.scala 66:30:@40155.4]
  assign _T_95185 = _T_95182[2]; // @[OneHot.scala 66:30:@40156.4]
  assign _T_95186 = _T_95182[3]; // @[OneHot.scala 66:30:@40157.4]
  assign _T_95187 = _T_95182[4]; // @[OneHot.scala 66:30:@40158.4]
  assign _T_95188 = _T_95182[5]; // @[OneHot.scala 66:30:@40159.4]
  assign _T_95189 = _T_95182[6]; // @[OneHot.scala 66:30:@40160.4]
  assign _T_95190 = _T_95182[7]; // @[OneHot.scala 66:30:@40161.4]
  assign _T_95191 = _T_95182[8]; // @[OneHot.scala 66:30:@40162.4]
  assign _T_95192 = _T_95182[9]; // @[OneHot.scala 66:30:@40163.4]
  assign _T_95193 = _T_95182[10]; // @[OneHot.scala 66:30:@40164.4]
  assign _T_95194 = _T_95182[11]; // @[OneHot.scala 66:30:@40165.4]
  assign _T_95195 = _T_95182[12]; // @[OneHot.scala 66:30:@40166.4]
  assign _T_95196 = _T_95182[13]; // @[OneHot.scala 66:30:@40167.4]
  assign _T_95197 = _T_95182[14]; // @[OneHot.scala 66:30:@40168.4]
  assign _T_95198 = _T_95182[15]; // @[OneHot.scala 66:30:@40169.4]
  assign _T_95239 = _T_94349 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40187.4]
  assign _T_95240 = _T_94346 ? 16'h4000 : _T_95239; // @[Mux.scala 31:69:@40188.4]
  assign _T_95241 = _T_94343 ? 16'h2000 : _T_95240; // @[Mux.scala 31:69:@40189.4]
  assign _T_95242 = _T_94340 ? 16'h1000 : _T_95241; // @[Mux.scala 31:69:@40190.4]
  assign _T_95243 = _T_94337 ? 16'h800 : _T_95242; // @[Mux.scala 31:69:@40191.4]
  assign _T_95244 = _T_94334 ? 16'h400 : _T_95243; // @[Mux.scala 31:69:@40192.4]
  assign _T_95245 = _T_94331 ? 16'h200 : _T_95244; // @[Mux.scala 31:69:@40193.4]
  assign _T_95246 = _T_94328 ? 16'h100 : _T_95245; // @[Mux.scala 31:69:@40194.4]
  assign _T_95247 = _T_94325 ? 16'h80 : _T_95246; // @[Mux.scala 31:69:@40195.4]
  assign _T_95248 = _T_94322 ? 16'h40 : _T_95247; // @[Mux.scala 31:69:@40196.4]
  assign _T_95249 = _T_94319 ? 16'h20 : _T_95248; // @[Mux.scala 31:69:@40197.4]
  assign _T_95250 = _T_94364 ? 16'h10 : _T_95249; // @[Mux.scala 31:69:@40198.4]
  assign _T_95251 = _T_94361 ? 16'h8 : _T_95250; // @[Mux.scala 31:69:@40199.4]
  assign _T_95252 = _T_94358 ? 16'h4 : _T_95251; // @[Mux.scala 31:69:@40200.4]
  assign _T_95253 = _T_94355 ? 16'h2 : _T_95252; // @[Mux.scala 31:69:@40201.4]
  assign _T_95254 = _T_94352 ? 16'h1 : _T_95253; // @[Mux.scala 31:69:@40202.4]
  assign _T_95255 = _T_95254[0]; // @[OneHot.scala 66:30:@40203.4]
  assign _T_95256 = _T_95254[1]; // @[OneHot.scala 66:30:@40204.4]
  assign _T_95257 = _T_95254[2]; // @[OneHot.scala 66:30:@40205.4]
  assign _T_95258 = _T_95254[3]; // @[OneHot.scala 66:30:@40206.4]
  assign _T_95259 = _T_95254[4]; // @[OneHot.scala 66:30:@40207.4]
  assign _T_95260 = _T_95254[5]; // @[OneHot.scala 66:30:@40208.4]
  assign _T_95261 = _T_95254[6]; // @[OneHot.scala 66:30:@40209.4]
  assign _T_95262 = _T_95254[7]; // @[OneHot.scala 66:30:@40210.4]
  assign _T_95263 = _T_95254[8]; // @[OneHot.scala 66:30:@40211.4]
  assign _T_95264 = _T_95254[9]; // @[OneHot.scala 66:30:@40212.4]
  assign _T_95265 = _T_95254[10]; // @[OneHot.scala 66:30:@40213.4]
  assign _T_95266 = _T_95254[11]; // @[OneHot.scala 66:30:@40214.4]
  assign _T_95267 = _T_95254[12]; // @[OneHot.scala 66:30:@40215.4]
  assign _T_95268 = _T_95254[13]; // @[OneHot.scala 66:30:@40216.4]
  assign _T_95269 = _T_95254[14]; // @[OneHot.scala 66:30:@40217.4]
  assign _T_95270 = _T_95254[15]; // @[OneHot.scala 66:30:@40218.4]
  assign _T_95311 = _T_94352 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40236.4]
  assign _T_95312 = _T_94349 ? 16'h4000 : _T_95311; // @[Mux.scala 31:69:@40237.4]
  assign _T_95313 = _T_94346 ? 16'h2000 : _T_95312; // @[Mux.scala 31:69:@40238.4]
  assign _T_95314 = _T_94343 ? 16'h1000 : _T_95313; // @[Mux.scala 31:69:@40239.4]
  assign _T_95315 = _T_94340 ? 16'h800 : _T_95314; // @[Mux.scala 31:69:@40240.4]
  assign _T_95316 = _T_94337 ? 16'h400 : _T_95315; // @[Mux.scala 31:69:@40241.4]
  assign _T_95317 = _T_94334 ? 16'h200 : _T_95316; // @[Mux.scala 31:69:@40242.4]
  assign _T_95318 = _T_94331 ? 16'h100 : _T_95317; // @[Mux.scala 31:69:@40243.4]
  assign _T_95319 = _T_94328 ? 16'h80 : _T_95318; // @[Mux.scala 31:69:@40244.4]
  assign _T_95320 = _T_94325 ? 16'h40 : _T_95319; // @[Mux.scala 31:69:@40245.4]
  assign _T_95321 = _T_94322 ? 16'h20 : _T_95320; // @[Mux.scala 31:69:@40246.4]
  assign _T_95322 = _T_94319 ? 16'h10 : _T_95321; // @[Mux.scala 31:69:@40247.4]
  assign _T_95323 = _T_94364 ? 16'h8 : _T_95322; // @[Mux.scala 31:69:@40248.4]
  assign _T_95324 = _T_94361 ? 16'h4 : _T_95323; // @[Mux.scala 31:69:@40249.4]
  assign _T_95325 = _T_94358 ? 16'h2 : _T_95324; // @[Mux.scala 31:69:@40250.4]
  assign _T_95326 = _T_94355 ? 16'h1 : _T_95325; // @[Mux.scala 31:69:@40251.4]
  assign _T_95327 = _T_95326[0]; // @[OneHot.scala 66:30:@40252.4]
  assign _T_95328 = _T_95326[1]; // @[OneHot.scala 66:30:@40253.4]
  assign _T_95329 = _T_95326[2]; // @[OneHot.scala 66:30:@40254.4]
  assign _T_95330 = _T_95326[3]; // @[OneHot.scala 66:30:@40255.4]
  assign _T_95331 = _T_95326[4]; // @[OneHot.scala 66:30:@40256.4]
  assign _T_95332 = _T_95326[5]; // @[OneHot.scala 66:30:@40257.4]
  assign _T_95333 = _T_95326[6]; // @[OneHot.scala 66:30:@40258.4]
  assign _T_95334 = _T_95326[7]; // @[OneHot.scala 66:30:@40259.4]
  assign _T_95335 = _T_95326[8]; // @[OneHot.scala 66:30:@40260.4]
  assign _T_95336 = _T_95326[9]; // @[OneHot.scala 66:30:@40261.4]
  assign _T_95337 = _T_95326[10]; // @[OneHot.scala 66:30:@40262.4]
  assign _T_95338 = _T_95326[11]; // @[OneHot.scala 66:30:@40263.4]
  assign _T_95339 = _T_95326[12]; // @[OneHot.scala 66:30:@40264.4]
  assign _T_95340 = _T_95326[13]; // @[OneHot.scala 66:30:@40265.4]
  assign _T_95341 = _T_95326[14]; // @[OneHot.scala 66:30:@40266.4]
  assign _T_95342 = _T_95326[15]; // @[OneHot.scala 66:30:@40267.4]
  assign _T_95383 = _T_94355 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40285.4]
  assign _T_95384 = _T_94352 ? 16'h4000 : _T_95383; // @[Mux.scala 31:69:@40286.4]
  assign _T_95385 = _T_94349 ? 16'h2000 : _T_95384; // @[Mux.scala 31:69:@40287.4]
  assign _T_95386 = _T_94346 ? 16'h1000 : _T_95385; // @[Mux.scala 31:69:@40288.4]
  assign _T_95387 = _T_94343 ? 16'h800 : _T_95386; // @[Mux.scala 31:69:@40289.4]
  assign _T_95388 = _T_94340 ? 16'h400 : _T_95387; // @[Mux.scala 31:69:@40290.4]
  assign _T_95389 = _T_94337 ? 16'h200 : _T_95388; // @[Mux.scala 31:69:@40291.4]
  assign _T_95390 = _T_94334 ? 16'h100 : _T_95389; // @[Mux.scala 31:69:@40292.4]
  assign _T_95391 = _T_94331 ? 16'h80 : _T_95390; // @[Mux.scala 31:69:@40293.4]
  assign _T_95392 = _T_94328 ? 16'h40 : _T_95391; // @[Mux.scala 31:69:@40294.4]
  assign _T_95393 = _T_94325 ? 16'h20 : _T_95392; // @[Mux.scala 31:69:@40295.4]
  assign _T_95394 = _T_94322 ? 16'h10 : _T_95393; // @[Mux.scala 31:69:@40296.4]
  assign _T_95395 = _T_94319 ? 16'h8 : _T_95394; // @[Mux.scala 31:69:@40297.4]
  assign _T_95396 = _T_94364 ? 16'h4 : _T_95395; // @[Mux.scala 31:69:@40298.4]
  assign _T_95397 = _T_94361 ? 16'h2 : _T_95396; // @[Mux.scala 31:69:@40299.4]
  assign _T_95398 = _T_94358 ? 16'h1 : _T_95397; // @[Mux.scala 31:69:@40300.4]
  assign _T_95399 = _T_95398[0]; // @[OneHot.scala 66:30:@40301.4]
  assign _T_95400 = _T_95398[1]; // @[OneHot.scala 66:30:@40302.4]
  assign _T_95401 = _T_95398[2]; // @[OneHot.scala 66:30:@40303.4]
  assign _T_95402 = _T_95398[3]; // @[OneHot.scala 66:30:@40304.4]
  assign _T_95403 = _T_95398[4]; // @[OneHot.scala 66:30:@40305.4]
  assign _T_95404 = _T_95398[5]; // @[OneHot.scala 66:30:@40306.4]
  assign _T_95405 = _T_95398[6]; // @[OneHot.scala 66:30:@40307.4]
  assign _T_95406 = _T_95398[7]; // @[OneHot.scala 66:30:@40308.4]
  assign _T_95407 = _T_95398[8]; // @[OneHot.scala 66:30:@40309.4]
  assign _T_95408 = _T_95398[9]; // @[OneHot.scala 66:30:@40310.4]
  assign _T_95409 = _T_95398[10]; // @[OneHot.scala 66:30:@40311.4]
  assign _T_95410 = _T_95398[11]; // @[OneHot.scala 66:30:@40312.4]
  assign _T_95411 = _T_95398[12]; // @[OneHot.scala 66:30:@40313.4]
  assign _T_95412 = _T_95398[13]; // @[OneHot.scala 66:30:@40314.4]
  assign _T_95413 = _T_95398[14]; // @[OneHot.scala 66:30:@40315.4]
  assign _T_95414 = _T_95398[15]; // @[OneHot.scala 66:30:@40316.4]
  assign _T_95455 = _T_94358 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40334.4]
  assign _T_95456 = _T_94355 ? 16'h4000 : _T_95455; // @[Mux.scala 31:69:@40335.4]
  assign _T_95457 = _T_94352 ? 16'h2000 : _T_95456; // @[Mux.scala 31:69:@40336.4]
  assign _T_95458 = _T_94349 ? 16'h1000 : _T_95457; // @[Mux.scala 31:69:@40337.4]
  assign _T_95459 = _T_94346 ? 16'h800 : _T_95458; // @[Mux.scala 31:69:@40338.4]
  assign _T_95460 = _T_94343 ? 16'h400 : _T_95459; // @[Mux.scala 31:69:@40339.4]
  assign _T_95461 = _T_94340 ? 16'h200 : _T_95460; // @[Mux.scala 31:69:@40340.4]
  assign _T_95462 = _T_94337 ? 16'h100 : _T_95461; // @[Mux.scala 31:69:@40341.4]
  assign _T_95463 = _T_94334 ? 16'h80 : _T_95462; // @[Mux.scala 31:69:@40342.4]
  assign _T_95464 = _T_94331 ? 16'h40 : _T_95463; // @[Mux.scala 31:69:@40343.4]
  assign _T_95465 = _T_94328 ? 16'h20 : _T_95464; // @[Mux.scala 31:69:@40344.4]
  assign _T_95466 = _T_94325 ? 16'h10 : _T_95465; // @[Mux.scala 31:69:@40345.4]
  assign _T_95467 = _T_94322 ? 16'h8 : _T_95466; // @[Mux.scala 31:69:@40346.4]
  assign _T_95468 = _T_94319 ? 16'h4 : _T_95467; // @[Mux.scala 31:69:@40347.4]
  assign _T_95469 = _T_94364 ? 16'h2 : _T_95468; // @[Mux.scala 31:69:@40348.4]
  assign _T_95470 = _T_94361 ? 16'h1 : _T_95469; // @[Mux.scala 31:69:@40349.4]
  assign _T_95471 = _T_95470[0]; // @[OneHot.scala 66:30:@40350.4]
  assign _T_95472 = _T_95470[1]; // @[OneHot.scala 66:30:@40351.4]
  assign _T_95473 = _T_95470[2]; // @[OneHot.scala 66:30:@40352.4]
  assign _T_95474 = _T_95470[3]; // @[OneHot.scala 66:30:@40353.4]
  assign _T_95475 = _T_95470[4]; // @[OneHot.scala 66:30:@40354.4]
  assign _T_95476 = _T_95470[5]; // @[OneHot.scala 66:30:@40355.4]
  assign _T_95477 = _T_95470[6]; // @[OneHot.scala 66:30:@40356.4]
  assign _T_95478 = _T_95470[7]; // @[OneHot.scala 66:30:@40357.4]
  assign _T_95479 = _T_95470[8]; // @[OneHot.scala 66:30:@40358.4]
  assign _T_95480 = _T_95470[9]; // @[OneHot.scala 66:30:@40359.4]
  assign _T_95481 = _T_95470[10]; // @[OneHot.scala 66:30:@40360.4]
  assign _T_95482 = _T_95470[11]; // @[OneHot.scala 66:30:@40361.4]
  assign _T_95483 = _T_95470[12]; // @[OneHot.scala 66:30:@40362.4]
  assign _T_95484 = _T_95470[13]; // @[OneHot.scala 66:30:@40363.4]
  assign _T_95485 = _T_95470[14]; // @[OneHot.scala 66:30:@40364.4]
  assign _T_95486 = _T_95470[15]; // @[OneHot.scala 66:30:@40365.4]
  assign _T_95527 = _T_94361 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40383.4]
  assign _T_95528 = _T_94358 ? 16'h4000 : _T_95527; // @[Mux.scala 31:69:@40384.4]
  assign _T_95529 = _T_94355 ? 16'h2000 : _T_95528; // @[Mux.scala 31:69:@40385.4]
  assign _T_95530 = _T_94352 ? 16'h1000 : _T_95529; // @[Mux.scala 31:69:@40386.4]
  assign _T_95531 = _T_94349 ? 16'h800 : _T_95530; // @[Mux.scala 31:69:@40387.4]
  assign _T_95532 = _T_94346 ? 16'h400 : _T_95531; // @[Mux.scala 31:69:@40388.4]
  assign _T_95533 = _T_94343 ? 16'h200 : _T_95532; // @[Mux.scala 31:69:@40389.4]
  assign _T_95534 = _T_94340 ? 16'h100 : _T_95533; // @[Mux.scala 31:69:@40390.4]
  assign _T_95535 = _T_94337 ? 16'h80 : _T_95534; // @[Mux.scala 31:69:@40391.4]
  assign _T_95536 = _T_94334 ? 16'h40 : _T_95535; // @[Mux.scala 31:69:@40392.4]
  assign _T_95537 = _T_94331 ? 16'h20 : _T_95536; // @[Mux.scala 31:69:@40393.4]
  assign _T_95538 = _T_94328 ? 16'h10 : _T_95537; // @[Mux.scala 31:69:@40394.4]
  assign _T_95539 = _T_94325 ? 16'h8 : _T_95538; // @[Mux.scala 31:69:@40395.4]
  assign _T_95540 = _T_94322 ? 16'h4 : _T_95539; // @[Mux.scala 31:69:@40396.4]
  assign _T_95541 = _T_94319 ? 16'h2 : _T_95540; // @[Mux.scala 31:69:@40397.4]
  assign _T_95542 = _T_94364 ? 16'h1 : _T_95541; // @[Mux.scala 31:69:@40398.4]
  assign _T_95543 = _T_95542[0]; // @[OneHot.scala 66:30:@40399.4]
  assign _T_95544 = _T_95542[1]; // @[OneHot.scala 66:30:@40400.4]
  assign _T_95545 = _T_95542[2]; // @[OneHot.scala 66:30:@40401.4]
  assign _T_95546 = _T_95542[3]; // @[OneHot.scala 66:30:@40402.4]
  assign _T_95547 = _T_95542[4]; // @[OneHot.scala 66:30:@40403.4]
  assign _T_95548 = _T_95542[5]; // @[OneHot.scala 66:30:@40404.4]
  assign _T_95549 = _T_95542[6]; // @[OneHot.scala 66:30:@40405.4]
  assign _T_95550 = _T_95542[7]; // @[OneHot.scala 66:30:@40406.4]
  assign _T_95551 = _T_95542[8]; // @[OneHot.scala 66:30:@40407.4]
  assign _T_95552 = _T_95542[9]; // @[OneHot.scala 66:30:@40408.4]
  assign _T_95553 = _T_95542[10]; // @[OneHot.scala 66:30:@40409.4]
  assign _T_95554 = _T_95542[11]; // @[OneHot.scala 66:30:@40410.4]
  assign _T_95555 = _T_95542[12]; // @[OneHot.scala 66:30:@40411.4]
  assign _T_95556 = _T_95542[13]; // @[OneHot.scala 66:30:@40412.4]
  assign _T_95557 = _T_95542[14]; // @[OneHot.scala 66:30:@40413.4]
  assign _T_95558 = _T_95542[15]; // @[OneHot.scala 66:30:@40414.4]
  assign _T_95623 = {_T_94470,_T_94469,_T_94468,_T_94467,_T_94466,_T_94465,_T_94464,_T_94463}; // @[Mux.scala 19:72:@40438.4]
  assign _T_95631 = {_T_94478,_T_94477,_T_94476,_T_94475,_T_94474,_T_94473,_T_94472,_T_94471,_T_95623}; // @[Mux.scala 19:72:@40446.4]
  assign _T_95633 = _T_90406 ? _T_95631 : 16'h0; // @[Mux.scala 19:72:@40447.4]
  assign _T_95640 = {_T_94541,_T_94540,_T_94539,_T_94538,_T_94537,_T_94536,_T_94535,_T_94550}; // @[Mux.scala 19:72:@40454.4]
  assign _T_95648 = {_T_94549,_T_94548,_T_94547,_T_94546,_T_94545,_T_94544,_T_94543,_T_94542,_T_95640}; // @[Mux.scala 19:72:@40462.4]
  assign _T_95650 = _T_90407 ? _T_95648 : 16'h0; // @[Mux.scala 19:72:@40463.4]
  assign _T_95657 = {_T_94612,_T_94611,_T_94610,_T_94609,_T_94608,_T_94607,_T_94622,_T_94621}; // @[Mux.scala 19:72:@40470.4]
  assign _T_95665 = {_T_94620,_T_94619,_T_94618,_T_94617,_T_94616,_T_94615,_T_94614,_T_94613,_T_95657}; // @[Mux.scala 19:72:@40478.4]
  assign _T_95667 = _T_90408 ? _T_95665 : 16'h0; // @[Mux.scala 19:72:@40479.4]
  assign _T_95674 = {_T_94683,_T_94682,_T_94681,_T_94680,_T_94679,_T_94694,_T_94693,_T_94692}; // @[Mux.scala 19:72:@40486.4]
  assign _T_95682 = {_T_94691,_T_94690,_T_94689,_T_94688,_T_94687,_T_94686,_T_94685,_T_94684,_T_95674}; // @[Mux.scala 19:72:@40494.4]
  assign _T_95684 = _T_90409 ? _T_95682 : 16'h0; // @[Mux.scala 19:72:@40495.4]
  assign _T_95691 = {_T_94754,_T_94753,_T_94752,_T_94751,_T_94766,_T_94765,_T_94764,_T_94763}; // @[Mux.scala 19:72:@40502.4]
  assign _T_95699 = {_T_94762,_T_94761,_T_94760,_T_94759,_T_94758,_T_94757,_T_94756,_T_94755,_T_95691}; // @[Mux.scala 19:72:@40510.4]
  assign _T_95701 = _T_90410 ? _T_95699 : 16'h0; // @[Mux.scala 19:72:@40511.4]
  assign _T_95708 = {_T_94825,_T_94824,_T_94823,_T_94838,_T_94837,_T_94836,_T_94835,_T_94834}; // @[Mux.scala 19:72:@40518.4]
  assign _T_95716 = {_T_94833,_T_94832,_T_94831,_T_94830,_T_94829,_T_94828,_T_94827,_T_94826,_T_95708}; // @[Mux.scala 19:72:@40526.4]
  assign _T_95718 = _T_90411 ? _T_95716 : 16'h0; // @[Mux.scala 19:72:@40527.4]
  assign _T_95725 = {_T_94896,_T_94895,_T_94910,_T_94909,_T_94908,_T_94907,_T_94906,_T_94905}; // @[Mux.scala 19:72:@40534.4]
  assign _T_95733 = {_T_94904,_T_94903,_T_94902,_T_94901,_T_94900,_T_94899,_T_94898,_T_94897,_T_95725}; // @[Mux.scala 19:72:@40542.4]
  assign _T_95735 = _T_90412 ? _T_95733 : 16'h0; // @[Mux.scala 19:72:@40543.4]
  assign _T_95742 = {_T_94967,_T_94982,_T_94981,_T_94980,_T_94979,_T_94978,_T_94977,_T_94976}; // @[Mux.scala 19:72:@40550.4]
  assign _T_95750 = {_T_94975,_T_94974,_T_94973,_T_94972,_T_94971,_T_94970,_T_94969,_T_94968,_T_95742}; // @[Mux.scala 19:72:@40558.4]
  assign _T_95752 = _T_90413 ? _T_95750 : 16'h0; // @[Mux.scala 19:72:@40559.4]
  assign _T_95759 = {_T_95054,_T_95053,_T_95052,_T_95051,_T_95050,_T_95049,_T_95048,_T_95047}; // @[Mux.scala 19:72:@40566.4]
  assign _T_95767 = {_T_95046,_T_95045,_T_95044,_T_95043,_T_95042,_T_95041,_T_95040,_T_95039,_T_95759}; // @[Mux.scala 19:72:@40574.4]
  assign _T_95769 = _T_90414 ? _T_95767 : 16'h0; // @[Mux.scala 19:72:@40575.4]
  assign _T_95776 = {_T_95125,_T_95124,_T_95123,_T_95122,_T_95121,_T_95120,_T_95119,_T_95118}; // @[Mux.scala 19:72:@40582.4]
  assign _T_95784 = {_T_95117,_T_95116,_T_95115,_T_95114,_T_95113,_T_95112,_T_95111,_T_95126,_T_95776}; // @[Mux.scala 19:72:@40590.4]
  assign _T_95786 = _T_90415 ? _T_95784 : 16'h0; // @[Mux.scala 19:72:@40591.4]
  assign _T_95793 = {_T_95196,_T_95195,_T_95194,_T_95193,_T_95192,_T_95191,_T_95190,_T_95189}; // @[Mux.scala 19:72:@40598.4]
  assign _T_95801 = {_T_95188,_T_95187,_T_95186,_T_95185,_T_95184,_T_95183,_T_95198,_T_95197,_T_95793}; // @[Mux.scala 19:72:@40606.4]
  assign _T_95803 = _T_90416 ? _T_95801 : 16'h0; // @[Mux.scala 19:72:@40607.4]
  assign _T_95810 = {_T_95267,_T_95266,_T_95265,_T_95264,_T_95263,_T_95262,_T_95261,_T_95260}; // @[Mux.scala 19:72:@40614.4]
  assign _T_95818 = {_T_95259,_T_95258,_T_95257,_T_95256,_T_95255,_T_95270,_T_95269,_T_95268,_T_95810}; // @[Mux.scala 19:72:@40622.4]
  assign _T_95820 = _T_90417 ? _T_95818 : 16'h0; // @[Mux.scala 19:72:@40623.4]
  assign _T_95827 = {_T_95338,_T_95337,_T_95336,_T_95335,_T_95334,_T_95333,_T_95332,_T_95331}; // @[Mux.scala 19:72:@40630.4]
  assign _T_95835 = {_T_95330,_T_95329,_T_95328,_T_95327,_T_95342,_T_95341,_T_95340,_T_95339,_T_95827}; // @[Mux.scala 19:72:@40638.4]
  assign _T_95837 = _T_90418 ? _T_95835 : 16'h0; // @[Mux.scala 19:72:@40639.4]
  assign _T_95844 = {_T_95409,_T_95408,_T_95407,_T_95406,_T_95405,_T_95404,_T_95403,_T_95402}; // @[Mux.scala 19:72:@40646.4]
  assign _T_95852 = {_T_95401,_T_95400,_T_95399,_T_95414,_T_95413,_T_95412,_T_95411,_T_95410,_T_95844}; // @[Mux.scala 19:72:@40654.4]
  assign _T_95854 = _T_90419 ? _T_95852 : 16'h0; // @[Mux.scala 19:72:@40655.4]
  assign _T_95861 = {_T_95480,_T_95479,_T_95478,_T_95477,_T_95476,_T_95475,_T_95474,_T_95473}; // @[Mux.scala 19:72:@40662.4]
  assign _T_95869 = {_T_95472,_T_95471,_T_95486,_T_95485,_T_95484,_T_95483,_T_95482,_T_95481,_T_95861}; // @[Mux.scala 19:72:@40670.4]
  assign _T_95871 = _T_90420 ? _T_95869 : 16'h0; // @[Mux.scala 19:72:@40671.4]
  assign _T_95878 = {_T_95551,_T_95550,_T_95549,_T_95548,_T_95547,_T_95546,_T_95545,_T_95544}; // @[Mux.scala 19:72:@40678.4]
  assign _T_95886 = {_T_95543,_T_95558,_T_95557,_T_95556,_T_95555,_T_95554,_T_95553,_T_95552,_T_95878}; // @[Mux.scala 19:72:@40686.4]
  assign _T_95888 = _T_90421 ? _T_95886 : 16'h0; // @[Mux.scala 19:72:@40687.4]
  assign _T_95889 = _T_95633 | _T_95650; // @[Mux.scala 19:72:@40688.4]
  assign _T_95890 = _T_95889 | _T_95667; // @[Mux.scala 19:72:@40689.4]
  assign _T_95891 = _T_95890 | _T_95684; // @[Mux.scala 19:72:@40690.4]
  assign _T_95892 = _T_95891 | _T_95701; // @[Mux.scala 19:72:@40691.4]
  assign _T_95893 = _T_95892 | _T_95718; // @[Mux.scala 19:72:@40692.4]
  assign _T_95894 = _T_95893 | _T_95735; // @[Mux.scala 19:72:@40693.4]
  assign _T_95895 = _T_95894 | _T_95752; // @[Mux.scala 19:72:@40694.4]
  assign _T_95896 = _T_95895 | _T_95769; // @[Mux.scala 19:72:@40695.4]
  assign _T_95897 = _T_95896 | _T_95786; // @[Mux.scala 19:72:@40696.4]
  assign _T_95898 = _T_95897 | _T_95803; // @[Mux.scala 19:72:@40697.4]
  assign _T_95899 = _T_95898 | _T_95820; // @[Mux.scala 19:72:@40698.4]
  assign _T_95900 = _T_95899 | _T_95837; // @[Mux.scala 19:72:@40699.4]
  assign _T_95901 = _T_95900 | _T_95854; // @[Mux.scala 19:72:@40700.4]
  assign _T_95902 = _T_95901 | _T_95871; // @[Mux.scala 19:72:@40701.4]
  assign _T_95903 = _T_95902 | _T_95888; // @[Mux.scala 19:72:@40702.4]
  assign inputPriorityPorts_0_0 = _T_95903[0]; // @[Mux.scala 19:72:@40706.4]
  assign inputPriorityPorts_0_1 = _T_95903[1]; // @[Mux.scala 19:72:@40708.4]
  assign inputPriorityPorts_0_2 = _T_95903[2]; // @[Mux.scala 19:72:@40710.4]
  assign inputPriorityPorts_0_3 = _T_95903[3]; // @[Mux.scala 19:72:@40712.4]
  assign inputPriorityPorts_0_4 = _T_95903[4]; // @[Mux.scala 19:72:@40714.4]
  assign inputPriorityPorts_0_5 = _T_95903[5]; // @[Mux.scala 19:72:@40716.4]
  assign inputPriorityPorts_0_6 = _T_95903[6]; // @[Mux.scala 19:72:@40718.4]
  assign inputPriorityPorts_0_7 = _T_95903[7]; // @[Mux.scala 19:72:@40720.4]
  assign inputPriorityPorts_0_8 = _T_95903[8]; // @[Mux.scala 19:72:@40722.4]
  assign inputPriorityPorts_0_9 = _T_95903[9]; // @[Mux.scala 19:72:@40724.4]
  assign inputPriorityPorts_0_10 = _T_95903[10]; // @[Mux.scala 19:72:@40726.4]
  assign inputPriorityPorts_0_11 = _T_95903[11]; // @[Mux.scala 19:72:@40728.4]
  assign inputPriorityPorts_0_12 = _T_95903[12]; // @[Mux.scala 19:72:@40730.4]
  assign inputPriorityPorts_0_13 = _T_95903[13]; // @[Mux.scala 19:72:@40732.4]
  assign inputPriorityPorts_0_14 = _T_95903[14]; // @[Mux.scala 19:72:@40734.4]
  assign inputPriorityPorts_0_15 = _T_95903[15]; // @[Mux.scala 19:72:@40736.4]
  assign _T_96105 = entriesPorts_0_15 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40790.4]
  assign _T_96106 = entriesPorts_0_14 ? 16'h4000 : _T_96105; // @[Mux.scala 31:69:@40791.4]
  assign _T_96107 = entriesPorts_0_13 ? 16'h2000 : _T_96106; // @[Mux.scala 31:69:@40792.4]
  assign _T_96108 = entriesPorts_0_12 ? 16'h1000 : _T_96107; // @[Mux.scala 31:69:@40793.4]
  assign _T_96109 = entriesPorts_0_11 ? 16'h800 : _T_96108; // @[Mux.scala 31:69:@40794.4]
  assign _T_96110 = entriesPorts_0_10 ? 16'h400 : _T_96109; // @[Mux.scala 31:69:@40795.4]
  assign _T_96111 = entriesPorts_0_9 ? 16'h200 : _T_96110; // @[Mux.scala 31:69:@40796.4]
  assign _T_96112 = entriesPorts_0_8 ? 16'h100 : _T_96111; // @[Mux.scala 31:69:@40797.4]
  assign _T_96113 = entriesPorts_0_7 ? 16'h80 : _T_96112; // @[Mux.scala 31:69:@40798.4]
  assign _T_96114 = entriesPorts_0_6 ? 16'h40 : _T_96113; // @[Mux.scala 31:69:@40799.4]
  assign _T_96115 = entriesPorts_0_5 ? 16'h20 : _T_96114; // @[Mux.scala 31:69:@40800.4]
  assign _T_96116 = entriesPorts_0_4 ? 16'h10 : _T_96115; // @[Mux.scala 31:69:@40801.4]
  assign _T_96117 = entriesPorts_0_3 ? 16'h8 : _T_96116; // @[Mux.scala 31:69:@40802.4]
  assign _T_96118 = entriesPorts_0_2 ? 16'h4 : _T_96117; // @[Mux.scala 31:69:@40803.4]
  assign _T_96119 = entriesPorts_0_1 ? 16'h2 : _T_96118; // @[Mux.scala 31:69:@40804.4]
  assign _T_96120 = entriesPorts_0_0 ? 16'h1 : _T_96119; // @[Mux.scala 31:69:@40805.4]
  assign _T_96121 = _T_96120[0]; // @[OneHot.scala 66:30:@40806.4]
  assign _T_96122 = _T_96120[1]; // @[OneHot.scala 66:30:@40807.4]
  assign _T_96123 = _T_96120[2]; // @[OneHot.scala 66:30:@40808.4]
  assign _T_96124 = _T_96120[3]; // @[OneHot.scala 66:30:@40809.4]
  assign _T_96125 = _T_96120[4]; // @[OneHot.scala 66:30:@40810.4]
  assign _T_96126 = _T_96120[5]; // @[OneHot.scala 66:30:@40811.4]
  assign _T_96127 = _T_96120[6]; // @[OneHot.scala 66:30:@40812.4]
  assign _T_96128 = _T_96120[7]; // @[OneHot.scala 66:30:@40813.4]
  assign _T_96129 = _T_96120[8]; // @[OneHot.scala 66:30:@40814.4]
  assign _T_96130 = _T_96120[9]; // @[OneHot.scala 66:30:@40815.4]
  assign _T_96131 = _T_96120[10]; // @[OneHot.scala 66:30:@40816.4]
  assign _T_96132 = _T_96120[11]; // @[OneHot.scala 66:30:@40817.4]
  assign _T_96133 = _T_96120[12]; // @[OneHot.scala 66:30:@40818.4]
  assign _T_96134 = _T_96120[13]; // @[OneHot.scala 66:30:@40819.4]
  assign _T_96135 = _T_96120[14]; // @[OneHot.scala 66:30:@40820.4]
  assign _T_96136 = _T_96120[15]; // @[OneHot.scala 66:30:@40821.4]
  assign _T_96177 = entriesPorts_0_0 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40839.4]
  assign _T_96178 = entriesPorts_0_15 ? 16'h4000 : _T_96177; // @[Mux.scala 31:69:@40840.4]
  assign _T_96179 = entriesPorts_0_14 ? 16'h2000 : _T_96178; // @[Mux.scala 31:69:@40841.4]
  assign _T_96180 = entriesPorts_0_13 ? 16'h1000 : _T_96179; // @[Mux.scala 31:69:@40842.4]
  assign _T_96181 = entriesPorts_0_12 ? 16'h800 : _T_96180; // @[Mux.scala 31:69:@40843.4]
  assign _T_96182 = entriesPorts_0_11 ? 16'h400 : _T_96181; // @[Mux.scala 31:69:@40844.4]
  assign _T_96183 = entriesPorts_0_10 ? 16'h200 : _T_96182; // @[Mux.scala 31:69:@40845.4]
  assign _T_96184 = entriesPorts_0_9 ? 16'h100 : _T_96183; // @[Mux.scala 31:69:@40846.4]
  assign _T_96185 = entriesPorts_0_8 ? 16'h80 : _T_96184; // @[Mux.scala 31:69:@40847.4]
  assign _T_96186 = entriesPorts_0_7 ? 16'h40 : _T_96185; // @[Mux.scala 31:69:@40848.4]
  assign _T_96187 = entriesPorts_0_6 ? 16'h20 : _T_96186; // @[Mux.scala 31:69:@40849.4]
  assign _T_96188 = entriesPorts_0_5 ? 16'h10 : _T_96187; // @[Mux.scala 31:69:@40850.4]
  assign _T_96189 = entriesPorts_0_4 ? 16'h8 : _T_96188; // @[Mux.scala 31:69:@40851.4]
  assign _T_96190 = entriesPorts_0_3 ? 16'h4 : _T_96189; // @[Mux.scala 31:69:@40852.4]
  assign _T_96191 = entriesPorts_0_2 ? 16'h2 : _T_96190; // @[Mux.scala 31:69:@40853.4]
  assign _T_96192 = entriesPorts_0_1 ? 16'h1 : _T_96191; // @[Mux.scala 31:69:@40854.4]
  assign _T_96193 = _T_96192[0]; // @[OneHot.scala 66:30:@40855.4]
  assign _T_96194 = _T_96192[1]; // @[OneHot.scala 66:30:@40856.4]
  assign _T_96195 = _T_96192[2]; // @[OneHot.scala 66:30:@40857.4]
  assign _T_96196 = _T_96192[3]; // @[OneHot.scala 66:30:@40858.4]
  assign _T_96197 = _T_96192[4]; // @[OneHot.scala 66:30:@40859.4]
  assign _T_96198 = _T_96192[5]; // @[OneHot.scala 66:30:@40860.4]
  assign _T_96199 = _T_96192[6]; // @[OneHot.scala 66:30:@40861.4]
  assign _T_96200 = _T_96192[7]; // @[OneHot.scala 66:30:@40862.4]
  assign _T_96201 = _T_96192[8]; // @[OneHot.scala 66:30:@40863.4]
  assign _T_96202 = _T_96192[9]; // @[OneHot.scala 66:30:@40864.4]
  assign _T_96203 = _T_96192[10]; // @[OneHot.scala 66:30:@40865.4]
  assign _T_96204 = _T_96192[11]; // @[OneHot.scala 66:30:@40866.4]
  assign _T_96205 = _T_96192[12]; // @[OneHot.scala 66:30:@40867.4]
  assign _T_96206 = _T_96192[13]; // @[OneHot.scala 66:30:@40868.4]
  assign _T_96207 = _T_96192[14]; // @[OneHot.scala 66:30:@40869.4]
  assign _T_96208 = _T_96192[15]; // @[OneHot.scala 66:30:@40870.4]
  assign _T_96249 = entriesPorts_0_1 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40888.4]
  assign _T_96250 = entriesPorts_0_0 ? 16'h4000 : _T_96249; // @[Mux.scala 31:69:@40889.4]
  assign _T_96251 = entriesPorts_0_15 ? 16'h2000 : _T_96250; // @[Mux.scala 31:69:@40890.4]
  assign _T_96252 = entriesPorts_0_14 ? 16'h1000 : _T_96251; // @[Mux.scala 31:69:@40891.4]
  assign _T_96253 = entriesPorts_0_13 ? 16'h800 : _T_96252; // @[Mux.scala 31:69:@40892.4]
  assign _T_96254 = entriesPorts_0_12 ? 16'h400 : _T_96253; // @[Mux.scala 31:69:@40893.4]
  assign _T_96255 = entriesPorts_0_11 ? 16'h200 : _T_96254; // @[Mux.scala 31:69:@40894.4]
  assign _T_96256 = entriesPorts_0_10 ? 16'h100 : _T_96255; // @[Mux.scala 31:69:@40895.4]
  assign _T_96257 = entriesPorts_0_9 ? 16'h80 : _T_96256; // @[Mux.scala 31:69:@40896.4]
  assign _T_96258 = entriesPorts_0_8 ? 16'h40 : _T_96257; // @[Mux.scala 31:69:@40897.4]
  assign _T_96259 = entriesPorts_0_7 ? 16'h20 : _T_96258; // @[Mux.scala 31:69:@40898.4]
  assign _T_96260 = entriesPorts_0_6 ? 16'h10 : _T_96259; // @[Mux.scala 31:69:@40899.4]
  assign _T_96261 = entriesPorts_0_5 ? 16'h8 : _T_96260; // @[Mux.scala 31:69:@40900.4]
  assign _T_96262 = entriesPorts_0_4 ? 16'h4 : _T_96261; // @[Mux.scala 31:69:@40901.4]
  assign _T_96263 = entriesPorts_0_3 ? 16'h2 : _T_96262; // @[Mux.scala 31:69:@40902.4]
  assign _T_96264 = entriesPorts_0_2 ? 16'h1 : _T_96263; // @[Mux.scala 31:69:@40903.4]
  assign _T_96265 = _T_96264[0]; // @[OneHot.scala 66:30:@40904.4]
  assign _T_96266 = _T_96264[1]; // @[OneHot.scala 66:30:@40905.4]
  assign _T_96267 = _T_96264[2]; // @[OneHot.scala 66:30:@40906.4]
  assign _T_96268 = _T_96264[3]; // @[OneHot.scala 66:30:@40907.4]
  assign _T_96269 = _T_96264[4]; // @[OneHot.scala 66:30:@40908.4]
  assign _T_96270 = _T_96264[5]; // @[OneHot.scala 66:30:@40909.4]
  assign _T_96271 = _T_96264[6]; // @[OneHot.scala 66:30:@40910.4]
  assign _T_96272 = _T_96264[7]; // @[OneHot.scala 66:30:@40911.4]
  assign _T_96273 = _T_96264[8]; // @[OneHot.scala 66:30:@40912.4]
  assign _T_96274 = _T_96264[9]; // @[OneHot.scala 66:30:@40913.4]
  assign _T_96275 = _T_96264[10]; // @[OneHot.scala 66:30:@40914.4]
  assign _T_96276 = _T_96264[11]; // @[OneHot.scala 66:30:@40915.4]
  assign _T_96277 = _T_96264[12]; // @[OneHot.scala 66:30:@40916.4]
  assign _T_96278 = _T_96264[13]; // @[OneHot.scala 66:30:@40917.4]
  assign _T_96279 = _T_96264[14]; // @[OneHot.scala 66:30:@40918.4]
  assign _T_96280 = _T_96264[15]; // @[OneHot.scala 66:30:@40919.4]
  assign _T_96321 = entriesPorts_0_2 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40937.4]
  assign _T_96322 = entriesPorts_0_1 ? 16'h4000 : _T_96321; // @[Mux.scala 31:69:@40938.4]
  assign _T_96323 = entriesPorts_0_0 ? 16'h2000 : _T_96322; // @[Mux.scala 31:69:@40939.4]
  assign _T_96324 = entriesPorts_0_15 ? 16'h1000 : _T_96323; // @[Mux.scala 31:69:@40940.4]
  assign _T_96325 = entriesPorts_0_14 ? 16'h800 : _T_96324; // @[Mux.scala 31:69:@40941.4]
  assign _T_96326 = entriesPorts_0_13 ? 16'h400 : _T_96325; // @[Mux.scala 31:69:@40942.4]
  assign _T_96327 = entriesPorts_0_12 ? 16'h200 : _T_96326; // @[Mux.scala 31:69:@40943.4]
  assign _T_96328 = entriesPorts_0_11 ? 16'h100 : _T_96327; // @[Mux.scala 31:69:@40944.4]
  assign _T_96329 = entriesPorts_0_10 ? 16'h80 : _T_96328; // @[Mux.scala 31:69:@40945.4]
  assign _T_96330 = entriesPorts_0_9 ? 16'h40 : _T_96329; // @[Mux.scala 31:69:@40946.4]
  assign _T_96331 = entriesPorts_0_8 ? 16'h20 : _T_96330; // @[Mux.scala 31:69:@40947.4]
  assign _T_96332 = entriesPorts_0_7 ? 16'h10 : _T_96331; // @[Mux.scala 31:69:@40948.4]
  assign _T_96333 = entriesPorts_0_6 ? 16'h8 : _T_96332; // @[Mux.scala 31:69:@40949.4]
  assign _T_96334 = entriesPorts_0_5 ? 16'h4 : _T_96333; // @[Mux.scala 31:69:@40950.4]
  assign _T_96335 = entriesPorts_0_4 ? 16'h2 : _T_96334; // @[Mux.scala 31:69:@40951.4]
  assign _T_96336 = entriesPorts_0_3 ? 16'h1 : _T_96335; // @[Mux.scala 31:69:@40952.4]
  assign _T_96337 = _T_96336[0]; // @[OneHot.scala 66:30:@40953.4]
  assign _T_96338 = _T_96336[1]; // @[OneHot.scala 66:30:@40954.4]
  assign _T_96339 = _T_96336[2]; // @[OneHot.scala 66:30:@40955.4]
  assign _T_96340 = _T_96336[3]; // @[OneHot.scala 66:30:@40956.4]
  assign _T_96341 = _T_96336[4]; // @[OneHot.scala 66:30:@40957.4]
  assign _T_96342 = _T_96336[5]; // @[OneHot.scala 66:30:@40958.4]
  assign _T_96343 = _T_96336[6]; // @[OneHot.scala 66:30:@40959.4]
  assign _T_96344 = _T_96336[7]; // @[OneHot.scala 66:30:@40960.4]
  assign _T_96345 = _T_96336[8]; // @[OneHot.scala 66:30:@40961.4]
  assign _T_96346 = _T_96336[9]; // @[OneHot.scala 66:30:@40962.4]
  assign _T_96347 = _T_96336[10]; // @[OneHot.scala 66:30:@40963.4]
  assign _T_96348 = _T_96336[11]; // @[OneHot.scala 66:30:@40964.4]
  assign _T_96349 = _T_96336[12]; // @[OneHot.scala 66:30:@40965.4]
  assign _T_96350 = _T_96336[13]; // @[OneHot.scala 66:30:@40966.4]
  assign _T_96351 = _T_96336[14]; // @[OneHot.scala 66:30:@40967.4]
  assign _T_96352 = _T_96336[15]; // @[OneHot.scala 66:30:@40968.4]
  assign _T_96393 = entriesPorts_0_3 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@40986.4]
  assign _T_96394 = entriesPorts_0_2 ? 16'h4000 : _T_96393; // @[Mux.scala 31:69:@40987.4]
  assign _T_96395 = entriesPorts_0_1 ? 16'h2000 : _T_96394; // @[Mux.scala 31:69:@40988.4]
  assign _T_96396 = entriesPorts_0_0 ? 16'h1000 : _T_96395; // @[Mux.scala 31:69:@40989.4]
  assign _T_96397 = entriesPorts_0_15 ? 16'h800 : _T_96396; // @[Mux.scala 31:69:@40990.4]
  assign _T_96398 = entriesPorts_0_14 ? 16'h400 : _T_96397; // @[Mux.scala 31:69:@40991.4]
  assign _T_96399 = entriesPorts_0_13 ? 16'h200 : _T_96398; // @[Mux.scala 31:69:@40992.4]
  assign _T_96400 = entriesPorts_0_12 ? 16'h100 : _T_96399; // @[Mux.scala 31:69:@40993.4]
  assign _T_96401 = entriesPorts_0_11 ? 16'h80 : _T_96400; // @[Mux.scala 31:69:@40994.4]
  assign _T_96402 = entriesPorts_0_10 ? 16'h40 : _T_96401; // @[Mux.scala 31:69:@40995.4]
  assign _T_96403 = entriesPorts_0_9 ? 16'h20 : _T_96402; // @[Mux.scala 31:69:@40996.4]
  assign _T_96404 = entriesPorts_0_8 ? 16'h10 : _T_96403; // @[Mux.scala 31:69:@40997.4]
  assign _T_96405 = entriesPorts_0_7 ? 16'h8 : _T_96404; // @[Mux.scala 31:69:@40998.4]
  assign _T_96406 = entriesPorts_0_6 ? 16'h4 : _T_96405; // @[Mux.scala 31:69:@40999.4]
  assign _T_96407 = entriesPorts_0_5 ? 16'h2 : _T_96406; // @[Mux.scala 31:69:@41000.4]
  assign _T_96408 = entriesPorts_0_4 ? 16'h1 : _T_96407; // @[Mux.scala 31:69:@41001.4]
  assign _T_96409 = _T_96408[0]; // @[OneHot.scala 66:30:@41002.4]
  assign _T_96410 = _T_96408[1]; // @[OneHot.scala 66:30:@41003.4]
  assign _T_96411 = _T_96408[2]; // @[OneHot.scala 66:30:@41004.4]
  assign _T_96412 = _T_96408[3]; // @[OneHot.scala 66:30:@41005.4]
  assign _T_96413 = _T_96408[4]; // @[OneHot.scala 66:30:@41006.4]
  assign _T_96414 = _T_96408[5]; // @[OneHot.scala 66:30:@41007.4]
  assign _T_96415 = _T_96408[6]; // @[OneHot.scala 66:30:@41008.4]
  assign _T_96416 = _T_96408[7]; // @[OneHot.scala 66:30:@41009.4]
  assign _T_96417 = _T_96408[8]; // @[OneHot.scala 66:30:@41010.4]
  assign _T_96418 = _T_96408[9]; // @[OneHot.scala 66:30:@41011.4]
  assign _T_96419 = _T_96408[10]; // @[OneHot.scala 66:30:@41012.4]
  assign _T_96420 = _T_96408[11]; // @[OneHot.scala 66:30:@41013.4]
  assign _T_96421 = _T_96408[12]; // @[OneHot.scala 66:30:@41014.4]
  assign _T_96422 = _T_96408[13]; // @[OneHot.scala 66:30:@41015.4]
  assign _T_96423 = _T_96408[14]; // @[OneHot.scala 66:30:@41016.4]
  assign _T_96424 = _T_96408[15]; // @[OneHot.scala 66:30:@41017.4]
  assign _T_96465 = entriesPorts_0_4 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41035.4]
  assign _T_96466 = entriesPorts_0_3 ? 16'h4000 : _T_96465; // @[Mux.scala 31:69:@41036.4]
  assign _T_96467 = entriesPorts_0_2 ? 16'h2000 : _T_96466; // @[Mux.scala 31:69:@41037.4]
  assign _T_96468 = entriesPorts_0_1 ? 16'h1000 : _T_96467; // @[Mux.scala 31:69:@41038.4]
  assign _T_96469 = entriesPorts_0_0 ? 16'h800 : _T_96468; // @[Mux.scala 31:69:@41039.4]
  assign _T_96470 = entriesPorts_0_15 ? 16'h400 : _T_96469; // @[Mux.scala 31:69:@41040.4]
  assign _T_96471 = entriesPorts_0_14 ? 16'h200 : _T_96470; // @[Mux.scala 31:69:@41041.4]
  assign _T_96472 = entriesPorts_0_13 ? 16'h100 : _T_96471; // @[Mux.scala 31:69:@41042.4]
  assign _T_96473 = entriesPorts_0_12 ? 16'h80 : _T_96472; // @[Mux.scala 31:69:@41043.4]
  assign _T_96474 = entriesPorts_0_11 ? 16'h40 : _T_96473; // @[Mux.scala 31:69:@41044.4]
  assign _T_96475 = entriesPorts_0_10 ? 16'h20 : _T_96474; // @[Mux.scala 31:69:@41045.4]
  assign _T_96476 = entriesPorts_0_9 ? 16'h10 : _T_96475; // @[Mux.scala 31:69:@41046.4]
  assign _T_96477 = entriesPorts_0_8 ? 16'h8 : _T_96476; // @[Mux.scala 31:69:@41047.4]
  assign _T_96478 = entriesPorts_0_7 ? 16'h4 : _T_96477; // @[Mux.scala 31:69:@41048.4]
  assign _T_96479 = entriesPorts_0_6 ? 16'h2 : _T_96478; // @[Mux.scala 31:69:@41049.4]
  assign _T_96480 = entriesPorts_0_5 ? 16'h1 : _T_96479; // @[Mux.scala 31:69:@41050.4]
  assign _T_96481 = _T_96480[0]; // @[OneHot.scala 66:30:@41051.4]
  assign _T_96482 = _T_96480[1]; // @[OneHot.scala 66:30:@41052.4]
  assign _T_96483 = _T_96480[2]; // @[OneHot.scala 66:30:@41053.4]
  assign _T_96484 = _T_96480[3]; // @[OneHot.scala 66:30:@41054.4]
  assign _T_96485 = _T_96480[4]; // @[OneHot.scala 66:30:@41055.4]
  assign _T_96486 = _T_96480[5]; // @[OneHot.scala 66:30:@41056.4]
  assign _T_96487 = _T_96480[6]; // @[OneHot.scala 66:30:@41057.4]
  assign _T_96488 = _T_96480[7]; // @[OneHot.scala 66:30:@41058.4]
  assign _T_96489 = _T_96480[8]; // @[OneHot.scala 66:30:@41059.4]
  assign _T_96490 = _T_96480[9]; // @[OneHot.scala 66:30:@41060.4]
  assign _T_96491 = _T_96480[10]; // @[OneHot.scala 66:30:@41061.4]
  assign _T_96492 = _T_96480[11]; // @[OneHot.scala 66:30:@41062.4]
  assign _T_96493 = _T_96480[12]; // @[OneHot.scala 66:30:@41063.4]
  assign _T_96494 = _T_96480[13]; // @[OneHot.scala 66:30:@41064.4]
  assign _T_96495 = _T_96480[14]; // @[OneHot.scala 66:30:@41065.4]
  assign _T_96496 = _T_96480[15]; // @[OneHot.scala 66:30:@41066.4]
  assign _T_96537 = entriesPorts_0_5 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41084.4]
  assign _T_96538 = entriesPorts_0_4 ? 16'h4000 : _T_96537; // @[Mux.scala 31:69:@41085.4]
  assign _T_96539 = entriesPorts_0_3 ? 16'h2000 : _T_96538; // @[Mux.scala 31:69:@41086.4]
  assign _T_96540 = entriesPorts_0_2 ? 16'h1000 : _T_96539; // @[Mux.scala 31:69:@41087.4]
  assign _T_96541 = entriesPorts_0_1 ? 16'h800 : _T_96540; // @[Mux.scala 31:69:@41088.4]
  assign _T_96542 = entriesPorts_0_0 ? 16'h400 : _T_96541; // @[Mux.scala 31:69:@41089.4]
  assign _T_96543 = entriesPorts_0_15 ? 16'h200 : _T_96542; // @[Mux.scala 31:69:@41090.4]
  assign _T_96544 = entriesPorts_0_14 ? 16'h100 : _T_96543; // @[Mux.scala 31:69:@41091.4]
  assign _T_96545 = entriesPorts_0_13 ? 16'h80 : _T_96544; // @[Mux.scala 31:69:@41092.4]
  assign _T_96546 = entriesPorts_0_12 ? 16'h40 : _T_96545; // @[Mux.scala 31:69:@41093.4]
  assign _T_96547 = entriesPorts_0_11 ? 16'h20 : _T_96546; // @[Mux.scala 31:69:@41094.4]
  assign _T_96548 = entriesPorts_0_10 ? 16'h10 : _T_96547; // @[Mux.scala 31:69:@41095.4]
  assign _T_96549 = entriesPorts_0_9 ? 16'h8 : _T_96548; // @[Mux.scala 31:69:@41096.4]
  assign _T_96550 = entriesPorts_0_8 ? 16'h4 : _T_96549; // @[Mux.scala 31:69:@41097.4]
  assign _T_96551 = entriesPorts_0_7 ? 16'h2 : _T_96550; // @[Mux.scala 31:69:@41098.4]
  assign _T_96552 = entriesPorts_0_6 ? 16'h1 : _T_96551; // @[Mux.scala 31:69:@41099.4]
  assign _T_96553 = _T_96552[0]; // @[OneHot.scala 66:30:@41100.4]
  assign _T_96554 = _T_96552[1]; // @[OneHot.scala 66:30:@41101.4]
  assign _T_96555 = _T_96552[2]; // @[OneHot.scala 66:30:@41102.4]
  assign _T_96556 = _T_96552[3]; // @[OneHot.scala 66:30:@41103.4]
  assign _T_96557 = _T_96552[4]; // @[OneHot.scala 66:30:@41104.4]
  assign _T_96558 = _T_96552[5]; // @[OneHot.scala 66:30:@41105.4]
  assign _T_96559 = _T_96552[6]; // @[OneHot.scala 66:30:@41106.4]
  assign _T_96560 = _T_96552[7]; // @[OneHot.scala 66:30:@41107.4]
  assign _T_96561 = _T_96552[8]; // @[OneHot.scala 66:30:@41108.4]
  assign _T_96562 = _T_96552[9]; // @[OneHot.scala 66:30:@41109.4]
  assign _T_96563 = _T_96552[10]; // @[OneHot.scala 66:30:@41110.4]
  assign _T_96564 = _T_96552[11]; // @[OneHot.scala 66:30:@41111.4]
  assign _T_96565 = _T_96552[12]; // @[OneHot.scala 66:30:@41112.4]
  assign _T_96566 = _T_96552[13]; // @[OneHot.scala 66:30:@41113.4]
  assign _T_96567 = _T_96552[14]; // @[OneHot.scala 66:30:@41114.4]
  assign _T_96568 = _T_96552[15]; // @[OneHot.scala 66:30:@41115.4]
  assign _T_96609 = entriesPorts_0_6 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41133.4]
  assign _T_96610 = entriesPorts_0_5 ? 16'h4000 : _T_96609; // @[Mux.scala 31:69:@41134.4]
  assign _T_96611 = entriesPorts_0_4 ? 16'h2000 : _T_96610; // @[Mux.scala 31:69:@41135.4]
  assign _T_96612 = entriesPorts_0_3 ? 16'h1000 : _T_96611; // @[Mux.scala 31:69:@41136.4]
  assign _T_96613 = entriesPorts_0_2 ? 16'h800 : _T_96612; // @[Mux.scala 31:69:@41137.4]
  assign _T_96614 = entriesPorts_0_1 ? 16'h400 : _T_96613; // @[Mux.scala 31:69:@41138.4]
  assign _T_96615 = entriesPorts_0_0 ? 16'h200 : _T_96614; // @[Mux.scala 31:69:@41139.4]
  assign _T_96616 = entriesPorts_0_15 ? 16'h100 : _T_96615; // @[Mux.scala 31:69:@41140.4]
  assign _T_96617 = entriesPorts_0_14 ? 16'h80 : _T_96616; // @[Mux.scala 31:69:@41141.4]
  assign _T_96618 = entriesPorts_0_13 ? 16'h40 : _T_96617; // @[Mux.scala 31:69:@41142.4]
  assign _T_96619 = entriesPorts_0_12 ? 16'h20 : _T_96618; // @[Mux.scala 31:69:@41143.4]
  assign _T_96620 = entriesPorts_0_11 ? 16'h10 : _T_96619; // @[Mux.scala 31:69:@41144.4]
  assign _T_96621 = entriesPorts_0_10 ? 16'h8 : _T_96620; // @[Mux.scala 31:69:@41145.4]
  assign _T_96622 = entriesPorts_0_9 ? 16'h4 : _T_96621; // @[Mux.scala 31:69:@41146.4]
  assign _T_96623 = entriesPorts_0_8 ? 16'h2 : _T_96622; // @[Mux.scala 31:69:@41147.4]
  assign _T_96624 = entriesPorts_0_7 ? 16'h1 : _T_96623; // @[Mux.scala 31:69:@41148.4]
  assign _T_96625 = _T_96624[0]; // @[OneHot.scala 66:30:@41149.4]
  assign _T_96626 = _T_96624[1]; // @[OneHot.scala 66:30:@41150.4]
  assign _T_96627 = _T_96624[2]; // @[OneHot.scala 66:30:@41151.4]
  assign _T_96628 = _T_96624[3]; // @[OneHot.scala 66:30:@41152.4]
  assign _T_96629 = _T_96624[4]; // @[OneHot.scala 66:30:@41153.4]
  assign _T_96630 = _T_96624[5]; // @[OneHot.scala 66:30:@41154.4]
  assign _T_96631 = _T_96624[6]; // @[OneHot.scala 66:30:@41155.4]
  assign _T_96632 = _T_96624[7]; // @[OneHot.scala 66:30:@41156.4]
  assign _T_96633 = _T_96624[8]; // @[OneHot.scala 66:30:@41157.4]
  assign _T_96634 = _T_96624[9]; // @[OneHot.scala 66:30:@41158.4]
  assign _T_96635 = _T_96624[10]; // @[OneHot.scala 66:30:@41159.4]
  assign _T_96636 = _T_96624[11]; // @[OneHot.scala 66:30:@41160.4]
  assign _T_96637 = _T_96624[12]; // @[OneHot.scala 66:30:@41161.4]
  assign _T_96638 = _T_96624[13]; // @[OneHot.scala 66:30:@41162.4]
  assign _T_96639 = _T_96624[14]; // @[OneHot.scala 66:30:@41163.4]
  assign _T_96640 = _T_96624[15]; // @[OneHot.scala 66:30:@41164.4]
  assign _T_96681 = entriesPorts_0_7 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41182.4]
  assign _T_96682 = entriesPorts_0_6 ? 16'h4000 : _T_96681; // @[Mux.scala 31:69:@41183.4]
  assign _T_96683 = entriesPorts_0_5 ? 16'h2000 : _T_96682; // @[Mux.scala 31:69:@41184.4]
  assign _T_96684 = entriesPorts_0_4 ? 16'h1000 : _T_96683; // @[Mux.scala 31:69:@41185.4]
  assign _T_96685 = entriesPorts_0_3 ? 16'h800 : _T_96684; // @[Mux.scala 31:69:@41186.4]
  assign _T_96686 = entriesPorts_0_2 ? 16'h400 : _T_96685; // @[Mux.scala 31:69:@41187.4]
  assign _T_96687 = entriesPorts_0_1 ? 16'h200 : _T_96686; // @[Mux.scala 31:69:@41188.4]
  assign _T_96688 = entriesPorts_0_0 ? 16'h100 : _T_96687; // @[Mux.scala 31:69:@41189.4]
  assign _T_96689 = entriesPorts_0_15 ? 16'h80 : _T_96688; // @[Mux.scala 31:69:@41190.4]
  assign _T_96690 = entriesPorts_0_14 ? 16'h40 : _T_96689; // @[Mux.scala 31:69:@41191.4]
  assign _T_96691 = entriesPorts_0_13 ? 16'h20 : _T_96690; // @[Mux.scala 31:69:@41192.4]
  assign _T_96692 = entriesPorts_0_12 ? 16'h10 : _T_96691; // @[Mux.scala 31:69:@41193.4]
  assign _T_96693 = entriesPorts_0_11 ? 16'h8 : _T_96692; // @[Mux.scala 31:69:@41194.4]
  assign _T_96694 = entriesPorts_0_10 ? 16'h4 : _T_96693; // @[Mux.scala 31:69:@41195.4]
  assign _T_96695 = entriesPorts_0_9 ? 16'h2 : _T_96694; // @[Mux.scala 31:69:@41196.4]
  assign _T_96696 = entriesPorts_0_8 ? 16'h1 : _T_96695; // @[Mux.scala 31:69:@41197.4]
  assign _T_96697 = _T_96696[0]; // @[OneHot.scala 66:30:@41198.4]
  assign _T_96698 = _T_96696[1]; // @[OneHot.scala 66:30:@41199.4]
  assign _T_96699 = _T_96696[2]; // @[OneHot.scala 66:30:@41200.4]
  assign _T_96700 = _T_96696[3]; // @[OneHot.scala 66:30:@41201.4]
  assign _T_96701 = _T_96696[4]; // @[OneHot.scala 66:30:@41202.4]
  assign _T_96702 = _T_96696[5]; // @[OneHot.scala 66:30:@41203.4]
  assign _T_96703 = _T_96696[6]; // @[OneHot.scala 66:30:@41204.4]
  assign _T_96704 = _T_96696[7]; // @[OneHot.scala 66:30:@41205.4]
  assign _T_96705 = _T_96696[8]; // @[OneHot.scala 66:30:@41206.4]
  assign _T_96706 = _T_96696[9]; // @[OneHot.scala 66:30:@41207.4]
  assign _T_96707 = _T_96696[10]; // @[OneHot.scala 66:30:@41208.4]
  assign _T_96708 = _T_96696[11]; // @[OneHot.scala 66:30:@41209.4]
  assign _T_96709 = _T_96696[12]; // @[OneHot.scala 66:30:@41210.4]
  assign _T_96710 = _T_96696[13]; // @[OneHot.scala 66:30:@41211.4]
  assign _T_96711 = _T_96696[14]; // @[OneHot.scala 66:30:@41212.4]
  assign _T_96712 = _T_96696[15]; // @[OneHot.scala 66:30:@41213.4]
  assign _T_96753 = entriesPorts_0_8 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41231.4]
  assign _T_96754 = entriesPorts_0_7 ? 16'h4000 : _T_96753; // @[Mux.scala 31:69:@41232.4]
  assign _T_96755 = entriesPorts_0_6 ? 16'h2000 : _T_96754; // @[Mux.scala 31:69:@41233.4]
  assign _T_96756 = entriesPorts_0_5 ? 16'h1000 : _T_96755; // @[Mux.scala 31:69:@41234.4]
  assign _T_96757 = entriesPorts_0_4 ? 16'h800 : _T_96756; // @[Mux.scala 31:69:@41235.4]
  assign _T_96758 = entriesPorts_0_3 ? 16'h400 : _T_96757; // @[Mux.scala 31:69:@41236.4]
  assign _T_96759 = entriesPorts_0_2 ? 16'h200 : _T_96758; // @[Mux.scala 31:69:@41237.4]
  assign _T_96760 = entriesPorts_0_1 ? 16'h100 : _T_96759; // @[Mux.scala 31:69:@41238.4]
  assign _T_96761 = entriesPorts_0_0 ? 16'h80 : _T_96760; // @[Mux.scala 31:69:@41239.4]
  assign _T_96762 = entriesPorts_0_15 ? 16'h40 : _T_96761; // @[Mux.scala 31:69:@41240.4]
  assign _T_96763 = entriesPorts_0_14 ? 16'h20 : _T_96762; // @[Mux.scala 31:69:@41241.4]
  assign _T_96764 = entriesPorts_0_13 ? 16'h10 : _T_96763; // @[Mux.scala 31:69:@41242.4]
  assign _T_96765 = entriesPorts_0_12 ? 16'h8 : _T_96764; // @[Mux.scala 31:69:@41243.4]
  assign _T_96766 = entriesPorts_0_11 ? 16'h4 : _T_96765; // @[Mux.scala 31:69:@41244.4]
  assign _T_96767 = entriesPorts_0_10 ? 16'h2 : _T_96766; // @[Mux.scala 31:69:@41245.4]
  assign _T_96768 = entriesPorts_0_9 ? 16'h1 : _T_96767; // @[Mux.scala 31:69:@41246.4]
  assign _T_96769 = _T_96768[0]; // @[OneHot.scala 66:30:@41247.4]
  assign _T_96770 = _T_96768[1]; // @[OneHot.scala 66:30:@41248.4]
  assign _T_96771 = _T_96768[2]; // @[OneHot.scala 66:30:@41249.4]
  assign _T_96772 = _T_96768[3]; // @[OneHot.scala 66:30:@41250.4]
  assign _T_96773 = _T_96768[4]; // @[OneHot.scala 66:30:@41251.4]
  assign _T_96774 = _T_96768[5]; // @[OneHot.scala 66:30:@41252.4]
  assign _T_96775 = _T_96768[6]; // @[OneHot.scala 66:30:@41253.4]
  assign _T_96776 = _T_96768[7]; // @[OneHot.scala 66:30:@41254.4]
  assign _T_96777 = _T_96768[8]; // @[OneHot.scala 66:30:@41255.4]
  assign _T_96778 = _T_96768[9]; // @[OneHot.scala 66:30:@41256.4]
  assign _T_96779 = _T_96768[10]; // @[OneHot.scala 66:30:@41257.4]
  assign _T_96780 = _T_96768[11]; // @[OneHot.scala 66:30:@41258.4]
  assign _T_96781 = _T_96768[12]; // @[OneHot.scala 66:30:@41259.4]
  assign _T_96782 = _T_96768[13]; // @[OneHot.scala 66:30:@41260.4]
  assign _T_96783 = _T_96768[14]; // @[OneHot.scala 66:30:@41261.4]
  assign _T_96784 = _T_96768[15]; // @[OneHot.scala 66:30:@41262.4]
  assign _T_96825 = entriesPorts_0_9 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41280.4]
  assign _T_96826 = entriesPorts_0_8 ? 16'h4000 : _T_96825; // @[Mux.scala 31:69:@41281.4]
  assign _T_96827 = entriesPorts_0_7 ? 16'h2000 : _T_96826; // @[Mux.scala 31:69:@41282.4]
  assign _T_96828 = entriesPorts_0_6 ? 16'h1000 : _T_96827; // @[Mux.scala 31:69:@41283.4]
  assign _T_96829 = entriesPorts_0_5 ? 16'h800 : _T_96828; // @[Mux.scala 31:69:@41284.4]
  assign _T_96830 = entriesPorts_0_4 ? 16'h400 : _T_96829; // @[Mux.scala 31:69:@41285.4]
  assign _T_96831 = entriesPorts_0_3 ? 16'h200 : _T_96830; // @[Mux.scala 31:69:@41286.4]
  assign _T_96832 = entriesPorts_0_2 ? 16'h100 : _T_96831; // @[Mux.scala 31:69:@41287.4]
  assign _T_96833 = entriesPorts_0_1 ? 16'h80 : _T_96832; // @[Mux.scala 31:69:@41288.4]
  assign _T_96834 = entriesPorts_0_0 ? 16'h40 : _T_96833; // @[Mux.scala 31:69:@41289.4]
  assign _T_96835 = entriesPorts_0_15 ? 16'h20 : _T_96834; // @[Mux.scala 31:69:@41290.4]
  assign _T_96836 = entriesPorts_0_14 ? 16'h10 : _T_96835; // @[Mux.scala 31:69:@41291.4]
  assign _T_96837 = entriesPorts_0_13 ? 16'h8 : _T_96836; // @[Mux.scala 31:69:@41292.4]
  assign _T_96838 = entriesPorts_0_12 ? 16'h4 : _T_96837; // @[Mux.scala 31:69:@41293.4]
  assign _T_96839 = entriesPorts_0_11 ? 16'h2 : _T_96838; // @[Mux.scala 31:69:@41294.4]
  assign _T_96840 = entriesPorts_0_10 ? 16'h1 : _T_96839; // @[Mux.scala 31:69:@41295.4]
  assign _T_96841 = _T_96840[0]; // @[OneHot.scala 66:30:@41296.4]
  assign _T_96842 = _T_96840[1]; // @[OneHot.scala 66:30:@41297.4]
  assign _T_96843 = _T_96840[2]; // @[OneHot.scala 66:30:@41298.4]
  assign _T_96844 = _T_96840[3]; // @[OneHot.scala 66:30:@41299.4]
  assign _T_96845 = _T_96840[4]; // @[OneHot.scala 66:30:@41300.4]
  assign _T_96846 = _T_96840[5]; // @[OneHot.scala 66:30:@41301.4]
  assign _T_96847 = _T_96840[6]; // @[OneHot.scala 66:30:@41302.4]
  assign _T_96848 = _T_96840[7]; // @[OneHot.scala 66:30:@41303.4]
  assign _T_96849 = _T_96840[8]; // @[OneHot.scala 66:30:@41304.4]
  assign _T_96850 = _T_96840[9]; // @[OneHot.scala 66:30:@41305.4]
  assign _T_96851 = _T_96840[10]; // @[OneHot.scala 66:30:@41306.4]
  assign _T_96852 = _T_96840[11]; // @[OneHot.scala 66:30:@41307.4]
  assign _T_96853 = _T_96840[12]; // @[OneHot.scala 66:30:@41308.4]
  assign _T_96854 = _T_96840[13]; // @[OneHot.scala 66:30:@41309.4]
  assign _T_96855 = _T_96840[14]; // @[OneHot.scala 66:30:@41310.4]
  assign _T_96856 = _T_96840[15]; // @[OneHot.scala 66:30:@41311.4]
  assign _T_96897 = entriesPorts_0_10 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41329.4]
  assign _T_96898 = entriesPorts_0_9 ? 16'h4000 : _T_96897; // @[Mux.scala 31:69:@41330.4]
  assign _T_96899 = entriesPorts_0_8 ? 16'h2000 : _T_96898; // @[Mux.scala 31:69:@41331.4]
  assign _T_96900 = entriesPorts_0_7 ? 16'h1000 : _T_96899; // @[Mux.scala 31:69:@41332.4]
  assign _T_96901 = entriesPorts_0_6 ? 16'h800 : _T_96900; // @[Mux.scala 31:69:@41333.4]
  assign _T_96902 = entriesPorts_0_5 ? 16'h400 : _T_96901; // @[Mux.scala 31:69:@41334.4]
  assign _T_96903 = entriesPorts_0_4 ? 16'h200 : _T_96902; // @[Mux.scala 31:69:@41335.4]
  assign _T_96904 = entriesPorts_0_3 ? 16'h100 : _T_96903; // @[Mux.scala 31:69:@41336.4]
  assign _T_96905 = entriesPorts_0_2 ? 16'h80 : _T_96904; // @[Mux.scala 31:69:@41337.4]
  assign _T_96906 = entriesPorts_0_1 ? 16'h40 : _T_96905; // @[Mux.scala 31:69:@41338.4]
  assign _T_96907 = entriesPorts_0_0 ? 16'h20 : _T_96906; // @[Mux.scala 31:69:@41339.4]
  assign _T_96908 = entriesPorts_0_15 ? 16'h10 : _T_96907; // @[Mux.scala 31:69:@41340.4]
  assign _T_96909 = entriesPorts_0_14 ? 16'h8 : _T_96908; // @[Mux.scala 31:69:@41341.4]
  assign _T_96910 = entriesPorts_0_13 ? 16'h4 : _T_96909; // @[Mux.scala 31:69:@41342.4]
  assign _T_96911 = entriesPorts_0_12 ? 16'h2 : _T_96910; // @[Mux.scala 31:69:@41343.4]
  assign _T_96912 = entriesPorts_0_11 ? 16'h1 : _T_96911; // @[Mux.scala 31:69:@41344.4]
  assign _T_96913 = _T_96912[0]; // @[OneHot.scala 66:30:@41345.4]
  assign _T_96914 = _T_96912[1]; // @[OneHot.scala 66:30:@41346.4]
  assign _T_96915 = _T_96912[2]; // @[OneHot.scala 66:30:@41347.4]
  assign _T_96916 = _T_96912[3]; // @[OneHot.scala 66:30:@41348.4]
  assign _T_96917 = _T_96912[4]; // @[OneHot.scala 66:30:@41349.4]
  assign _T_96918 = _T_96912[5]; // @[OneHot.scala 66:30:@41350.4]
  assign _T_96919 = _T_96912[6]; // @[OneHot.scala 66:30:@41351.4]
  assign _T_96920 = _T_96912[7]; // @[OneHot.scala 66:30:@41352.4]
  assign _T_96921 = _T_96912[8]; // @[OneHot.scala 66:30:@41353.4]
  assign _T_96922 = _T_96912[9]; // @[OneHot.scala 66:30:@41354.4]
  assign _T_96923 = _T_96912[10]; // @[OneHot.scala 66:30:@41355.4]
  assign _T_96924 = _T_96912[11]; // @[OneHot.scala 66:30:@41356.4]
  assign _T_96925 = _T_96912[12]; // @[OneHot.scala 66:30:@41357.4]
  assign _T_96926 = _T_96912[13]; // @[OneHot.scala 66:30:@41358.4]
  assign _T_96927 = _T_96912[14]; // @[OneHot.scala 66:30:@41359.4]
  assign _T_96928 = _T_96912[15]; // @[OneHot.scala 66:30:@41360.4]
  assign _T_96969 = entriesPorts_0_11 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41378.4]
  assign _T_96970 = entriesPorts_0_10 ? 16'h4000 : _T_96969; // @[Mux.scala 31:69:@41379.4]
  assign _T_96971 = entriesPorts_0_9 ? 16'h2000 : _T_96970; // @[Mux.scala 31:69:@41380.4]
  assign _T_96972 = entriesPorts_0_8 ? 16'h1000 : _T_96971; // @[Mux.scala 31:69:@41381.4]
  assign _T_96973 = entriesPorts_0_7 ? 16'h800 : _T_96972; // @[Mux.scala 31:69:@41382.4]
  assign _T_96974 = entriesPorts_0_6 ? 16'h400 : _T_96973; // @[Mux.scala 31:69:@41383.4]
  assign _T_96975 = entriesPorts_0_5 ? 16'h200 : _T_96974; // @[Mux.scala 31:69:@41384.4]
  assign _T_96976 = entriesPorts_0_4 ? 16'h100 : _T_96975; // @[Mux.scala 31:69:@41385.4]
  assign _T_96977 = entriesPorts_0_3 ? 16'h80 : _T_96976; // @[Mux.scala 31:69:@41386.4]
  assign _T_96978 = entriesPorts_0_2 ? 16'h40 : _T_96977; // @[Mux.scala 31:69:@41387.4]
  assign _T_96979 = entriesPorts_0_1 ? 16'h20 : _T_96978; // @[Mux.scala 31:69:@41388.4]
  assign _T_96980 = entriesPorts_0_0 ? 16'h10 : _T_96979; // @[Mux.scala 31:69:@41389.4]
  assign _T_96981 = entriesPorts_0_15 ? 16'h8 : _T_96980; // @[Mux.scala 31:69:@41390.4]
  assign _T_96982 = entriesPorts_0_14 ? 16'h4 : _T_96981; // @[Mux.scala 31:69:@41391.4]
  assign _T_96983 = entriesPorts_0_13 ? 16'h2 : _T_96982; // @[Mux.scala 31:69:@41392.4]
  assign _T_96984 = entriesPorts_0_12 ? 16'h1 : _T_96983; // @[Mux.scala 31:69:@41393.4]
  assign _T_96985 = _T_96984[0]; // @[OneHot.scala 66:30:@41394.4]
  assign _T_96986 = _T_96984[1]; // @[OneHot.scala 66:30:@41395.4]
  assign _T_96987 = _T_96984[2]; // @[OneHot.scala 66:30:@41396.4]
  assign _T_96988 = _T_96984[3]; // @[OneHot.scala 66:30:@41397.4]
  assign _T_96989 = _T_96984[4]; // @[OneHot.scala 66:30:@41398.4]
  assign _T_96990 = _T_96984[5]; // @[OneHot.scala 66:30:@41399.4]
  assign _T_96991 = _T_96984[6]; // @[OneHot.scala 66:30:@41400.4]
  assign _T_96992 = _T_96984[7]; // @[OneHot.scala 66:30:@41401.4]
  assign _T_96993 = _T_96984[8]; // @[OneHot.scala 66:30:@41402.4]
  assign _T_96994 = _T_96984[9]; // @[OneHot.scala 66:30:@41403.4]
  assign _T_96995 = _T_96984[10]; // @[OneHot.scala 66:30:@41404.4]
  assign _T_96996 = _T_96984[11]; // @[OneHot.scala 66:30:@41405.4]
  assign _T_96997 = _T_96984[12]; // @[OneHot.scala 66:30:@41406.4]
  assign _T_96998 = _T_96984[13]; // @[OneHot.scala 66:30:@41407.4]
  assign _T_96999 = _T_96984[14]; // @[OneHot.scala 66:30:@41408.4]
  assign _T_97000 = _T_96984[15]; // @[OneHot.scala 66:30:@41409.4]
  assign _T_97041 = entriesPorts_0_12 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41427.4]
  assign _T_97042 = entriesPorts_0_11 ? 16'h4000 : _T_97041; // @[Mux.scala 31:69:@41428.4]
  assign _T_97043 = entriesPorts_0_10 ? 16'h2000 : _T_97042; // @[Mux.scala 31:69:@41429.4]
  assign _T_97044 = entriesPorts_0_9 ? 16'h1000 : _T_97043; // @[Mux.scala 31:69:@41430.4]
  assign _T_97045 = entriesPorts_0_8 ? 16'h800 : _T_97044; // @[Mux.scala 31:69:@41431.4]
  assign _T_97046 = entriesPorts_0_7 ? 16'h400 : _T_97045; // @[Mux.scala 31:69:@41432.4]
  assign _T_97047 = entriesPorts_0_6 ? 16'h200 : _T_97046; // @[Mux.scala 31:69:@41433.4]
  assign _T_97048 = entriesPorts_0_5 ? 16'h100 : _T_97047; // @[Mux.scala 31:69:@41434.4]
  assign _T_97049 = entriesPorts_0_4 ? 16'h80 : _T_97048; // @[Mux.scala 31:69:@41435.4]
  assign _T_97050 = entriesPorts_0_3 ? 16'h40 : _T_97049; // @[Mux.scala 31:69:@41436.4]
  assign _T_97051 = entriesPorts_0_2 ? 16'h20 : _T_97050; // @[Mux.scala 31:69:@41437.4]
  assign _T_97052 = entriesPorts_0_1 ? 16'h10 : _T_97051; // @[Mux.scala 31:69:@41438.4]
  assign _T_97053 = entriesPorts_0_0 ? 16'h8 : _T_97052; // @[Mux.scala 31:69:@41439.4]
  assign _T_97054 = entriesPorts_0_15 ? 16'h4 : _T_97053; // @[Mux.scala 31:69:@41440.4]
  assign _T_97055 = entriesPorts_0_14 ? 16'h2 : _T_97054; // @[Mux.scala 31:69:@41441.4]
  assign _T_97056 = entriesPorts_0_13 ? 16'h1 : _T_97055; // @[Mux.scala 31:69:@41442.4]
  assign _T_97057 = _T_97056[0]; // @[OneHot.scala 66:30:@41443.4]
  assign _T_97058 = _T_97056[1]; // @[OneHot.scala 66:30:@41444.4]
  assign _T_97059 = _T_97056[2]; // @[OneHot.scala 66:30:@41445.4]
  assign _T_97060 = _T_97056[3]; // @[OneHot.scala 66:30:@41446.4]
  assign _T_97061 = _T_97056[4]; // @[OneHot.scala 66:30:@41447.4]
  assign _T_97062 = _T_97056[5]; // @[OneHot.scala 66:30:@41448.4]
  assign _T_97063 = _T_97056[6]; // @[OneHot.scala 66:30:@41449.4]
  assign _T_97064 = _T_97056[7]; // @[OneHot.scala 66:30:@41450.4]
  assign _T_97065 = _T_97056[8]; // @[OneHot.scala 66:30:@41451.4]
  assign _T_97066 = _T_97056[9]; // @[OneHot.scala 66:30:@41452.4]
  assign _T_97067 = _T_97056[10]; // @[OneHot.scala 66:30:@41453.4]
  assign _T_97068 = _T_97056[11]; // @[OneHot.scala 66:30:@41454.4]
  assign _T_97069 = _T_97056[12]; // @[OneHot.scala 66:30:@41455.4]
  assign _T_97070 = _T_97056[13]; // @[OneHot.scala 66:30:@41456.4]
  assign _T_97071 = _T_97056[14]; // @[OneHot.scala 66:30:@41457.4]
  assign _T_97072 = _T_97056[15]; // @[OneHot.scala 66:30:@41458.4]
  assign _T_97113 = entriesPorts_0_13 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41476.4]
  assign _T_97114 = entriesPorts_0_12 ? 16'h4000 : _T_97113; // @[Mux.scala 31:69:@41477.4]
  assign _T_97115 = entriesPorts_0_11 ? 16'h2000 : _T_97114; // @[Mux.scala 31:69:@41478.4]
  assign _T_97116 = entriesPorts_0_10 ? 16'h1000 : _T_97115; // @[Mux.scala 31:69:@41479.4]
  assign _T_97117 = entriesPorts_0_9 ? 16'h800 : _T_97116; // @[Mux.scala 31:69:@41480.4]
  assign _T_97118 = entriesPorts_0_8 ? 16'h400 : _T_97117; // @[Mux.scala 31:69:@41481.4]
  assign _T_97119 = entriesPorts_0_7 ? 16'h200 : _T_97118; // @[Mux.scala 31:69:@41482.4]
  assign _T_97120 = entriesPorts_0_6 ? 16'h100 : _T_97119; // @[Mux.scala 31:69:@41483.4]
  assign _T_97121 = entriesPorts_0_5 ? 16'h80 : _T_97120; // @[Mux.scala 31:69:@41484.4]
  assign _T_97122 = entriesPorts_0_4 ? 16'h40 : _T_97121; // @[Mux.scala 31:69:@41485.4]
  assign _T_97123 = entriesPorts_0_3 ? 16'h20 : _T_97122; // @[Mux.scala 31:69:@41486.4]
  assign _T_97124 = entriesPorts_0_2 ? 16'h10 : _T_97123; // @[Mux.scala 31:69:@41487.4]
  assign _T_97125 = entriesPorts_0_1 ? 16'h8 : _T_97124; // @[Mux.scala 31:69:@41488.4]
  assign _T_97126 = entriesPorts_0_0 ? 16'h4 : _T_97125; // @[Mux.scala 31:69:@41489.4]
  assign _T_97127 = entriesPorts_0_15 ? 16'h2 : _T_97126; // @[Mux.scala 31:69:@41490.4]
  assign _T_97128 = entriesPorts_0_14 ? 16'h1 : _T_97127; // @[Mux.scala 31:69:@41491.4]
  assign _T_97129 = _T_97128[0]; // @[OneHot.scala 66:30:@41492.4]
  assign _T_97130 = _T_97128[1]; // @[OneHot.scala 66:30:@41493.4]
  assign _T_97131 = _T_97128[2]; // @[OneHot.scala 66:30:@41494.4]
  assign _T_97132 = _T_97128[3]; // @[OneHot.scala 66:30:@41495.4]
  assign _T_97133 = _T_97128[4]; // @[OneHot.scala 66:30:@41496.4]
  assign _T_97134 = _T_97128[5]; // @[OneHot.scala 66:30:@41497.4]
  assign _T_97135 = _T_97128[6]; // @[OneHot.scala 66:30:@41498.4]
  assign _T_97136 = _T_97128[7]; // @[OneHot.scala 66:30:@41499.4]
  assign _T_97137 = _T_97128[8]; // @[OneHot.scala 66:30:@41500.4]
  assign _T_97138 = _T_97128[9]; // @[OneHot.scala 66:30:@41501.4]
  assign _T_97139 = _T_97128[10]; // @[OneHot.scala 66:30:@41502.4]
  assign _T_97140 = _T_97128[11]; // @[OneHot.scala 66:30:@41503.4]
  assign _T_97141 = _T_97128[12]; // @[OneHot.scala 66:30:@41504.4]
  assign _T_97142 = _T_97128[13]; // @[OneHot.scala 66:30:@41505.4]
  assign _T_97143 = _T_97128[14]; // @[OneHot.scala 66:30:@41506.4]
  assign _T_97144 = _T_97128[15]; // @[OneHot.scala 66:30:@41507.4]
  assign _T_97185 = entriesPorts_0_14 ? 16'h8000 : 16'h0; // @[Mux.scala 31:69:@41525.4]
  assign _T_97186 = entriesPorts_0_13 ? 16'h4000 : _T_97185; // @[Mux.scala 31:69:@41526.4]
  assign _T_97187 = entriesPorts_0_12 ? 16'h2000 : _T_97186; // @[Mux.scala 31:69:@41527.4]
  assign _T_97188 = entriesPorts_0_11 ? 16'h1000 : _T_97187; // @[Mux.scala 31:69:@41528.4]
  assign _T_97189 = entriesPorts_0_10 ? 16'h800 : _T_97188; // @[Mux.scala 31:69:@41529.4]
  assign _T_97190 = entriesPorts_0_9 ? 16'h400 : _T_97189; // @[Mux.scala 31:69:@41530.4]
  assign _T_97191 = entriesPorts_0_8 ? 16'h200 : _T_97190; // @[Mux.scala 31:69:@41531.4]
  assign _T_97192 = entriesPorts_0_7 ? 16'h100 : _T_97191; // @[Mux.scala 31:69:@41532.4]
  assign _T_97193 = entriesPorts_0_6 ? 16'h80 : _T_97192; // @[Mux.scala 31:69:@41533.4]
  assign _T_97194 = entriesPorts_0_5 ? 16'h40 : _T_97193; // @[Mux.scala 31:69:@41534.4]
  assign _T_97195 = entriesPorts_0_4 ? 16'h20 : _T_97194; // @[Mux.scala 31:69:@41535.4]
  assign _T_97196 = entriesPorts_0_3 ? 16'h10 : _T_97195; // @[Mux.scala 31:69:@41536.4]
  assign _T_97197 = entriesPorts_0_2 ? 16'h8 : _T_97196; // @[Mux.scala 31:69:@41537.4]
  assign _T_97198 = entriesPorts_0_1 ? 16'h4 : _T_97197; // @[Mux.scala 31:69:@41538.4]
  assign _T_97199 = entriesPorts_0_0 ? 16'h2 : _T_97198; // @[Mux.scala 31:69:@41539.4]
  assign _T_97200 = entriesPorts_0_15 ? 16'h1 : _T_97199; // @[Mux.scala 31:69:@41540.4]
  assign _T_97201 = _T_97200[0]; // @[OneHot.scala 66:30:@41541.4]
  assign _T_97202 = _T_97200[1]; // @[OneHot.scala 66:30:@41542.4]
  assign _T_97203 = _T_97200[2]; // @[OneHot.scala 66:30:@41543.4]
  assign _T_97204 = _T_97200[3]; // @[OneHot.scala 66:30:@41544.4]
  assign _T_97205 = _T_97200[4]; // @[OneHot.scala 66:30:@41545.4]
  assign _T_97206 = _T_97200[5]; // @[OneHot.scala 66:30:@41546.4]
  assign _T_97207 = _T_97200[6]; // @[OneHot.scala 66:30:@41547.4]
  assign _T_97208 = _T_97200[7]; // @[OneHot.scala 66:30:@41548.4]
  assign _T_97209 = _T_97200[8]; // @[OneHot.scala 66:30:@41549.4]
  assign _T_97210 = _T_97200[9]; // @[OneHot.scala 66:30:@41550.4]
  assign _T_97211 = _T_97200[10]; // @[OneHot.scala 66:30:@41551.4]
  assign _T_97212 = _T_97200[11]; // @[OneHot.scala 66:30:@41552.4]
  assign _T_97213 = _T_97200[12]; // @[OneHot.scala 66:30:@41553.4]
  assign _T_97214 = _T_97200[13]; // @[OneHot.scala 66:30:@41554.4]
  assign _T_97215 = _T_97200[14]; // @[OneHot.scala 66:30:@41555.4]
  assign _T_97216 = _T_97200[15]; // @[OneHot.scala 66:30:@41556.4]
  assign _T_97281 = {_T_96128,_T_96127,_T_96126,_T_96125,_T_96124,_T_96123,_T_96122,_T_96121}; // @[Mux.scala 19:72:@41580.4]
  assign _T_97289 = {_T_96136,_T_96135,_T_96134,_T_96133,_T_96132,_T_96131,_T_96130,_T_96129,_T_97281}; // @[Mux.scala 19:72:@41588.4]
  assign _T_97291 = _T_90406 ? _T_97289 : 16'h0; // @[Mux.scala 19:72:@41589.4]
  assign _T_97298 = {_T_96199,_T_96198,_T_96197,_T_96196,_T_96195,_T_96194,_T_96193,_T_96208}; // @[Mux.scala 19:72:@41596.4]
  assign _T_97306 = {_T_96207,_T_96206,_T_96205,_T_96204,_T_96203,_T_96202,_T_96201,_T_96200,_T_97298}; // @[Mux.scala 19:72:@41604.4]
  assign _T_97308 = _T_90407 ? _T_97306 : 16'h0; // @[Mux.scala 19:72:@41605.4]
  assign _T_97315 = {_T_96270,_T_96269,_T_96268,_T_96267,_T_96266,_T_96265,_T_96280,_T_96279}; // @[Mux.scala 19:72:@41612.4]
  assign _T_97323 = {_T_96278,_T_96277,_T_96276,_T_96275,_T_96274,_T_96273,_T_96272,_T_96271,_T_97315}; // @[Mux.scala 19:72:@41620.4]
  assign _T_97325 = _T_90408 ? _T_97323 : 16'h0; // @[Mux.scala 19:72:@41621.4]
  assign _T_97332 = {_T_96341,_T_96340,_T_96339,_T_96338,_T_96337,_T_96352,_T_96351,_T_96350}; // @[Mux.scala 19:72:@41628.4]
  assign _T_97340 = {_T_96349,_T_96348,_T_96347,_T_96346,_T_96345,_T_96344,_T_96343,_T_96342,_T_97332}; // @[Mux.scala 19:72:@41636.4]
  assign _T_97342 = _T_90409 ? _T_97340 : 16'h0; // @[Mux.scala 19:72:@41637.4]
  assign _T_97349 = {_T_96412,_T_96411,_T_96410,_T_96409,_T_96424,_T_96423,_T_96422,_T_96421}; // @[Mux.scala 19:72:@41644.4]
  assign _T_97357 = {_T_96420,_T_96419,_T_96418,_T_96417,_T_96416,_T_96415,_T_96414,_T_96413,_T_97349}; // @[Mux.scala 19:72:@41652.4]
  assign _T_97359 = _T_90410 ? _T_97357 : 16'h0; // @[Mux.scala 19:72:@41653.4]
  assign _T_97366 = {_T_96483,_T_96482,_T_96481,_T_96496,_T_96495,_T_96494,_T_96493,_T_96492}; // @[Mux.scala 19:72:@41660.4]
  assign _T_97374 = {_T_96491,_T_96490,_T_96489,_T_96488,_T_96487,_T_96486,_T_96485,_T_96484,_T_97366}; // @[Mux.scala 19:72:@41668.4]
  assign _T_97376 = _T_90411 ? _T_97374 : 16'h0; // @[Mux.scala 19:72:@41669.4]
  assign _T_97383 = {_T_96554,_T_96553,_T_96568,_T_96567,_T_96566,_T_96565,_T_96564,_T_96563}; // @[Mux.scala 19:72:@41676.4]
  assign _T_97391 = {_T_96562,_T_96561,_T_96560,_T_96559,_T_96558,_T_96557,_T_96556,_T_96555,_T_97383}; // @[Mux.scala 19:72:@41684.4]
  assign _T_97393 = _T_90412 ? _T_97391 : 16'h0; // @[Mux.scala 19:72:@41685.4]
  assign _T_97400 = {_T_96625,_T_96640,_T_96639,_T_96638,_T_96637,_T_96636,_T_96635,_T_96634}; // @[Mux.scala 19:72:@41692.4]
  assign _T_97408 = {_T_96633,_T_96632,_T_96631,_T_96630,_T_96629,_T_96628,_T_96627,_T_96626,_T_97400}; // @[Mux.scala 19:72:@41700.4]
  assign _T_97410 = _T_90413 ? _T_97408 : 16'h0; // @[Mux.scala 19:72:@41701.4]
  assign _T_97417 = {_T_96712,_T_96711,_T_96710,_T_96709,_T_96708,_T_96707,_T_96706,_T_96705}; // @[Mux.scala 19:72:@41708.4]
  assign _T_97425 = {_T_96704,_T_96703,_T_96702,_T_96701,_T_96700,_T_96699,_T_96698,_T_96697,_T_97417}; // @[Mux.scala 19:72:@41716.4]
  assign _T_97427 = _T_90414 ? _T_97425 : 16'h0; // @[Mux.scala 19:72:@41717.4]
  assign _T_97434 = {_T_96783,_T_96782,_T_96781,_T_96780,_T_96779,_T_96778,_T_96777,_T_96776}; // @[Mux.scala 19:72:@41724.4]
  assign _T_97442 = {_T_96775,_T_96774,_T_96773,_T_96772,_T_96771,_T_96770,_T_96769,_T_96784,_T_97434}; // @[Mux.scala 19:72:@41732.4]
  assign _T_97444 = _T_90415 ? _T_97442 : 16'h0; // @[Mux.scala 19:72:@41733.4]
  assign _T_97451 = {_T_96854,_T_96853,_T_96852,_T_96851,_T_96850,_T_96849,_T_96848,_T_96847}; // @[Mux.scala 19:72:@41740.4]
  assign _T_97459 = {_T_96846,_T_96845,_T_96844,_T_96843,_T_96842,_T_96841,_T_96856,_T_96855,_T_97451}; // @[Mux.scala 19:72:@41748.4]
  assign _T_97461 = _T_90416 ? _T_97459 : 16'h0; // @[Mux.scala 19:72:@41749.4]
  assign _T_97468 = {_T_96925,_T_96924,_T_96923,_T_96922,_T_96921,_T_96920,_T_96919,_T_96918}; // @[Mux.scala 19:72:@41756.4]
  assign _T_97476 = {_T_96917,_T_96916,_T_96915,_T_96914,_T_96913,_T_96928,_T_96927,_T_96926,_T_97468}; // @[Mux.scala 19:72:@41764.4]
  assign _T_97478 = _T_90417 ? _T_97476 : 16'h0; // @[Mux.scala 19:72:@41765.4]
  assign _T_97485 = {_T_96996,_T_96995,_T_96994,_T_96993,_T_96992,_T_96991,_T_96990,_T_96989}; // @[Mux.scala 19:72:@41772.4]
  assign _T_97493 = {_T_96988,_T_96987,_T_96986,_T_96985,_T_97000,_T_96999,_T_96998,_T_96997,_T_97485}; // @[Mux.scala 19:72:@41780.4]
  assign _T_97495 = _T_90418 ? _T_97493 : 16'h0; // @[Mux.scala 19:72:@41781.4]
  assign _T_97502 = {_T_97067,_T_97066,_T_97065,_T_97064,_T_97063,_T_97062,_T_97061,_T_97060}; // @[Mux.scala 19:72:@41788.4]
  assign _T_97510 = {_T_97059,_T_97058,_T_97057,_T_97072,_T_97071,_T_97070,_T_97069,_T_97068,_T_97502}; // @[Mux.scala 19:72:@41796.4]
  assign _T_97512 = _T_90419 ? _T_97510 : 16'h0; // @[Mux.scala 19:72:@41797.4]
  assign _T_97519 = {_T_97138,_T_97137,_T_97136,_T_97135,_T_97134,_T_97133,_T_97132,_T_97131}; // @[Mux.scala 19:72:@41804.4]
  assign _T_97527 = {_T_97130,_T_97129,_T_97144,_T_97143,_T_97142,_T_97141,_T_97140,_T_97139,_T_97519}; // @[Mux.scala 19:72:@41812.4]
  assign _T_97529 = _T_90420 ? _T_97527 : 16'h0; // @[Mux.scala 19:72:@41813.4]
  assign _T_97536 = {_T_97209,_T_97208,_T_97207,_T_97206,_T_97205,_T_97204,_T_97203,_T_97202}; // @[Mux.scala 19:72:@41820.4]
  assign _T_97544 = {_T_97201,_T_97216,_T_97215,_T_97214,_T_97213,_T_97212,_T_97211,_T_97210,_T_97536}; // @[Mux.scala 19:72:@41828.4]
  assign _T_97546 = _T_90421 ? _T_97544 : 16'h0; // @[Mux.scala 19:72:@41829.4]
  assign _T_97547 = _T_97291 | _T_97308; // @[Mux.scala 19:72:@41830.4]
  assign _T_97548 = _T_97547 | _T_97325; // @[Mux.scala 19:72:@41831.4]
  assign _T_97549 = _T_97548 | _T_97342; // @[Mux.scala 19:72:@41832.4]
  assign _T_97550 = _T_97549 | _T_97359; // @[Mux.scala 19:72:@41833.4]
  assign _T_97551 = _T_97550 | _T_97376; // @[Mux.scala 19:72:@41834.4]
  assign _T_97552 = _T_97551 | _T_97393; // @[Mux.scala 19:72:@41835.4]
  assign _T_97553 = _T_97552 | _T_97410; // @[Mux.scala 19:72:@41836.4]
  assign _T_97554 = _T_97553 | _T_97427; // @[Mux.scala 19:72:@41837.4]
  assign _T_97555 = _T_97554 | _T_97444; // @[Mux.scala 19:72:@41838.4]
  assign _T_97556 = _T_97555 | _T_97461; // @[Mux.scala 19:72:@41839.4]
  assign _T_97557 = _T_97556 | _T_97478; // @[Mux.scala 19:72:@41840.4]
  assign _T_97558 = _T_97557 | _T_97495; // @[Mux.scala 19:72:@41841.4]
  assign _T_97559 = _T_97558 | _T_97512; // @[Mux.scala 19:72:@41842.4]
  assign _T_97560 = _T_97559 | _T_97529; // @[Mux.scala 19:72:@41843.4]
  assign _T_97561 = _T_97560 | _T_97546; // @[Mux.scala 19:72:@41844.4]
  assign outputPriorityPorts_0_0 = _T_97561[0]; // @[Mux.scala 19:72:@41848.4]
  assign outputPriorityPorts_0_1 = _T_97561[1]; // @[Mux.scala 19:72:@41850.4]
  assign outputPriorityPorts_0_2 = _T_97561[2]; // @[Mux.scala 19:72:@41852.4]
  assign outputPriorityPorts_0_3 = _T_97561[3]; // @[Mux.scala 19:72:@41854.4]
  assign outputPriorityPorts_0_4 = _T_97561[4]; // @[Mux.scala 19:72:@41856.4]
  assign outputPriorityPorts_0_5 = _T_97561[5]; // @[Mux.scala 19:72:@41858.4]
  assign outputPriorityPorts_0_6 = _T_97561[6]; // @[Mux.scala 19:72:@41860.4]
  assign outputPriorityPorts_0_7 = _T_97561[7]; // @[Mux.scala 19:72:@41862.4]
  assign outputPriorityPorts_0_8 = _T_97561[8]; // @[Mux.scala 19:72:@41864.4]
  assign outputPriorityPorts_0_9 = _T_97561[9]; // @[Mux.scala 19:72:@41866.4]
  assign outputPriorityPorts_0_10 = _T_97561[10]; // @[Mux.scala 19:72:@41868.4]
  assign outputPriorityPorts_0_11 = _T_97561[11]; // @[Mux.scala 19:72:@41870.4]
  assign outputPriorityPorts_0_12 = _T_97561[12]; // @[Mux.scala 19:72:@41872.4]
  assign outputPriorityPorts_0_13 = _T_97561[13]; // @[Mux.scala 19:72:@41874.4]
  assign outputPriorityPorts_0_14 = _T_97561[14]; // @[Mux.scala 19:72:@41876.4]
  assign outputPriorityPorts_0_15 = _T_97561[15]; // @[Mux.scala 19:72:@41878.4]
  assign _T_97704 = inputPriorityPorts_0_0 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41900.6]
  assign _GEN_2128 = _T_97704 ? io_addrFromLoadPorts_0 : addrQ_0; // @[AxiLoadQueue.scala 316:36:@41904.6]
  assign _GEN_2129 = _T_97704 ? 1'h1 : addrKnown_0; // @[AxiLoadQueue.scala 316:36:@41904.6]
  assign _GEN_2130 = initBits_0 ? 1'h0 : _GEN_2129; // @[AxiLoadQueue.scala 310:34:@41896.4]
  assign _GEN_2131 = initBits_0 ? addrQ_0 : _GEN_2128; // @[AxiLoadQueue.scala 310:34:@41896.4]
  assign _T_97719 = inputPriorityPorts_0_1 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41913.6]
  assign _GEN_2132 = _T_97719 ? io_addrFromLoadPorts_0 : addrQ_1; // @[AxiLoadQueue.scala 316:36:@41917.6]
  assign _GEN_2133 = _T_97719 ? 1'h1 : addrKnown_1; // @[AxiLoadQueue.scala 316:36:@41917.6]
  assign _GEN_2134 = initBits_1 ? 1'h0 : _GEN_2133; // @[AxiLoadQueue.scala 310:34:@41909.4]
  assign _GEN_2135 = initBits_1 ? addrQ_1 : _GEN_2132; // @[AxiLoadQueue.scala 310:34:@41909.4]
  assign _T_97734 = inputPriorityPorts_0_2 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41926.6]
  assign _GEN_2136 = _T_97734 ? io_addrFromLoadPorts_0 : addrQ_2; // @[AxiLoadQueue.scala 316:36:@41930.6]
  assign _GEN_2137 = _T_97734 ? 1'h1 : addrKnown_2; // @[AxiLoadQueue.scala 316:36:@41930.6]
  assign _GEN_2138 = initBits_2 ? 1'h0 : _GEN_2137; // @[AxiLoadQueue.scala 310:34:@41922.4]
  assign _GEN_2139 = initBits_2 ? addrQ_2 : _GEN_2136; // @[AxiLoadQueue.scala 310:34:@41922.4]
  assign _T_97749 = inputPriorityPorts_0_3 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41939.6]
  assign _GEN_2140 = _T_97749 ? io_addrFromLoadPorts_0 : addrQ_3; // @[AxiLoadQueue.scala 316:36:@41943.6]
  assign _GEN_2141 = _T_97749 ? 1'h1 : addrKnown_3; // @[AxiLoadQueue.scala 316:36:@41943.6]
  assign _GEN_2142 = initBits_3 ? 1'h0 : _GEN_2141; // @[AxiLoadQueue.scala 310:34:@41935.4]
  assign _GEN_2143 = initBits_3 ? addrQ_3 : _GEN_2140; // @[AxiLoadQueue.scala 310:34:@41935.4]
  assign _T_97764 = inputPriorityPorts_0_4 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41952.6]
  assign _GEN_2144 = _T_97764 ? io_addrFromLoadPorts_0 : addrQ_4; // @[AxiLoadQueue.scala 316:36:@41956.6]
  assign _GEN_2145 = _T_97764 ? 1'h1 : addrKnown_4; // @[AxiLoadQueue.scala 316:36:@41956.6]
  assign _GEN_2146 = initBits_4 ? 1'h0 : _GEN_2145; // @[AxiLoadQueue.scala 310:34:@41948.4]
  assign _GEN_2147 = initBits_4 ? addrQ_4 : _GEN_2144; // @[AxiLoadQueue.scala 310:34:@41948.4]
  assign _T_97779 = inputPriorityPorts_0_5 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41965.6]
  assign _GEN_2148 = _T_97779 ? io_addrFromLoadPorts_0 : addrQ_5; // @[AxiLoadQueue.scala 316:36:@41969.6]
  assign _GEN_2149 = _T_97779 ? 1'h1 : addrKnown_5; // @[AxiLoadQueue.scala 316:36:@41969.6]
  assign _GEN_2150 = initBits_5 ? 1'h0 : _GEN_2149; // @[AxiLoadQueue.scala 310:34:@41961.4]
  assign _GEN_2151 = initBits_5 ? addrQ_5 : _GEN_2148; // @[AxiLoadQueue.scala 310:34:@41961.4]
  assign _T_97794 = inputPriorityPorts_0_6 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41978.6]
  assign _GEN_2152 = _T_97794 ? io_addrFromLoadPorts_0 : addrQ_6; // @[AxiLoadQueue.scala 316:36:@41982.6]
  assign _GEN_2153 = _T_97794 ? 1'h1 : addrKnown_6; // @[AxiLoadQueue.scala 316:36:@41982.6]
  assign _GEN_2154 = initBits_6 ? 1'h0 : _GEN_2153; // @[AxiLoadQueue.scala 310:34:@41974.4]
  assign _GEN_2155 = initBits_6 ? addrQ_6 : _GEN_2152; // @[AxiLoadQueue.scala 310:34:@41974.4]
  assign _T_97809 = inputPriorityPorts_0_7 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@41991.6]
  assign _GEN_2156 = _T_97809 ? io_addrFromLoadPorts_0 : addrQ_7; // @[AxiLoadQueue.scala 316:36:@41995.6]
  assign _GEN_2157 = _T_97809 ? 1'h1 : addrKnown_7; // @[AxiLoadQueue.scala 316:36:@41995.6]
  assign _GEN_2158 = initBits_7 ? 1'h0 : _GEN_2157; // @[AxiLoadQueue.scala 310:34:@41987.4]
  assign _GEN_2159 = initBits_7 ? addrQ_7 : _GEN_2156; // @[AxiLoadQueue.scala 310:34:@41987.4]
  assign _T_97824 = inputPriorityPorts_0_8 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42004.6]
  assign _GEN_2160 = _T_97824 ? io_addrFromLoadPorts_0 : addrQ_8; // @[AxiLoadQueue.scala 316:36:@42008.6]
  assign _GEN_2161 = _T_97824 ? 1'h1 : addrKnown_8; // @[AxiLoadQueue.scala 316:36:@42008.6]
  assign _GEN_2162 = initBits_8 ? 1'h0 : _GEN_2161; // @[AxiLoadQueue.scala 310:34:@42000.4]
  assign _GEN_2163 = initBits_8 ? addrQ_8 : _GEN_2160; // @[AxiLoadQueue.scala 310:34:@42000.4]
  assign _T_97839 = inputPriorityPorts_0_9 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42017.6]
  assign _GEN_2164 = _T_97839 ? io_addrFromLoadPorts_0 : addrQ_9; // @[AxiLoadQueue.scala 316:36:@42021.6]
  assign _GEN_2165 = _T_97839 ? 1'h1 : addrKnown_9; // @[AxiLoadQueue.scala 316:36:@42021.6]
  assign _GEN_2166 = initBits_9 ? 1'h0 : _GEN_2165; // @[AxiLoadQueue.scala 310:34:@42013.4]
  assign _GEN_2167 = initBits_9 ? addrQ_9 : _GEN_2164; // @[AxiLoadQueue.scala 310:34:@42013.4]
  assign _T_97854 = inputPriorityPorts_0_10 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42030.6]
  assign _GEN_2168 = _T_97854 ? io_addrFromLoadPorts_0 : addrQ_10; // @[AxiLoadQueue.scala 316:36:@42034.6]
  assign _GEN_2169 = _T_97854 ? 1'h1 : addrKnown_10; // @[AxiLoadQueue.scala 316:36:@42034.6]
  assign _GEN_2170 = initBits_10 ? 1'h0 : _GEN_2169; // @[AxiLoadQueue.scala 310:34:@42026.4]
  assign _GEN_2171 = initBits_10 ? addrQ_10 : _GEN_2168; // @[AxiLoadQueue.scala 310:34:@42026.4]
  assign _T_97869 = inputPriorityPorts_0_11 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42043.6]
  assign _GEN_2172 = _T_97869 ? io_addrFromLoadPorts_0 : addrQ_11; // @[AxiLoadQueue.scala 316:36:@42047.6]
  assign _GEN_2173 = _T_97869 ? 1'h1 : addrKnown_11; // @[AxiLoadQueue.scala 316:36:@42047.6]
  assign _GEN_2174 = initBits_11 ? 1'h0 : _GEN_2173; // @[AxiLoadQueue.scala 310:34:@42039.4]
  assign _GEN_2175 = initBits_11 ? addrQ_11 : _GEN_2172; // @[AxiLoadQueue.scala 310:34:@42039.4]
  assign _T_97884 = inputPriorityPorts_0_12 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42056.6]
  assign _GEN_2176 = _T_97884 ? io_addrFromLoadPorts_0 : addrQ_12; // @[AxiLoadQueue.scala 316:36:@42060.6]
  assign _GEN_2177 = _T_97884 ? 1'h1 : addrKnown_12; // @[AxiLoadQueue.scala 316:36:@42060.6]
  assign _GEN_2178 = initBits_12 ? 1'h0 : _GEN_2177; // @[AxiLoadQueue.scala 310:34:@42052.4]
  assign _GEN_2179 = initBits_12 ? addrQ_12 : _GEN_2176; // @[AxiLoadQueue.scala 310:34:@42052.4]
  assign _T_97899 = inputPriorityPorts_0_13 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42069.6]
  assign _GEN_2180 = _T_97899 ? io_addrFromLoadPorts_0 : addrQ_13; // @[AxiLoadQueue.scala 316:36:@42073.6]
  assign _GEN_2181 = _T_97899 ? 1'h1 : addrKnown_13; // @[AxiLoadQueue.scala 316:36:@42073.6]
  assign _GEN_2182 = initBits_13 ? 1'h0 : _GEN_2181; // @[AxiLoadQueue.scala 310:34:@42065.4]
  assign _GEN_2183 = initBits_13 ? addrQ_13 : _GEN_2180; // @[AxiLoadQueue.scala 310:34:@42065.4]
  assign _T_97914 = inputPriorityPorts_0_14 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42082.6]
  assign _GEN_2184 = _T_97914 ? io_addrFromLoadPorts_0 : addrQ_14; // @[AxiLoadQueue.scala 316:36:@42086.6]
  assign _GEN_2185 = _T_97914 ? 1'h1 : addrKnown_14; // @[AxiLoadQueue.scala 316:36:@42086.6]
  assign _GEN_2186 = initBits_14 ? 1'h0 : _GEN_2185; // @[AxiLoadQueue.scala 310:34:@42078.4]
  assign _GEN_2187 = initBits_14 ? addrQ_14 : _GEN_2184; // @[AxiLoadQueue.scala 310:34:@42078.4]
  assign _T_97929 = inputPriorityPorts_0_15 & io_loadAddrEnable_0; // @[AxiLoadQueue.scala 315:47:@42095.6]
  assign _GEN_2188 = _T_97929 ? io_addrFromLoadPorts_0 : addrQ_15; // @[AxiLoadQueue.scala 316:36:@42099.6]
  assign _GEN_2189 = _T_97929 ? 1'h1 : addrKnown_15; // @[AxiLoadQueue.scala 316:36:@42099.6]
  assign _GEN_2190 = initBits_15 ? 1'h0 : _GEN_2189; // @[AxiLoadQueue.scala 310:34:@42091.4]
  assign _GEN_2191 = initBits_15 ? addrQ_15 : _GEN_2188; // @[AxiLoadQueue.scala 310:34:@42091.4]
  assign _T_97964 = outputPriorityPorts_0_0 & dataKnown_0; // @[AxiLoadQueue.scala 328:108:@42105.4]
  assign _T_97966 = loadCompleted_0 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42106.4]
  assign _T_97967 = _T_97964 & _T_97966; // @[AxiLoadQueue.scala 329:31:@42107.4]
  assign loadCompleting_0 = _T_97967 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42108.4]
  assign _T_97978 = outputPriorityPorts_0_1 & dataKnown_1; // @[AxiLoadQueue.scala 328:108:@42113.4]
  assign _T_97980 = loadCompleted_1 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42114.4]
  assign _T_97981 = _T_97978 & _T_97980; // @[AxiLoadQueue.scala 329:31:@42115.4]
  assign loadCompleting_1 = _T_97981 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42116.4]
  assign _T_97992 = outputPriorityPorts_0_2 & dataKnown_2; // @[AxiLoadQueue.scala 328:108:@42121.4]
  assign _T_97994 = loadCompleted_2 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42122.4]
  assign _T_97995 = _T_97992 & _T_97994; // @[AxiLoadQueue.scala 329:31:@42123.4]
  assign loadCompleting_2 = _T_97995 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42124.4]
  assign _T_98006 = outputPriorityPorts_0_3 & dataKnown_3; // @[AxiLoadQueue.scala 328:108:@42129.4]
  assign _T_98008 = loadCompleted_3 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42130.4]
  assign _T_98009 = _T_98006 & _T_98008; // @[AxiLoadQueue.scala 329:31:@42131.4]
  assign loadCompleting_3 = _T_98009 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42132.4]
  assign _T_98020 = outputPriorityPorts_0_4 & dataKnown_4; // @[AxiLoadQueue.scala 328:108:@42137.4]
  assign _T_98022 = loadCompleted_4 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42138.4]
  assign _T_98023 = _T_98020 & _T_98022; // @[AxiLoadQueue.scala 329:31:@42139.4]
  assign loadCompleting_4 = _T_98023 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42140.4]
  assign _T_98034 = outputPriorityPorts_0_5 & dataKnown_5; // @[AxiLoadQueue.scala 328:108:@42145.4]
  assign _T_98036 = loadCompleted_5 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42146.4]
  assign _T_98037 = _T_98034 & _T_98036; // @[AxiLoadQueue.scala 329:31:@42147.4]
  assign loadCompleting_5 = _T_98037 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42148.4]
  assign _T_98048 = outputPriorityPorts_0_6 & dataKnown_6; // @[AxiLoadQueue.scala 328:108:@42153.4]
  assign _T_98050 = loadCompleted_6 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42154.4]
  assign _T_98051 = _T_98048 & _T_98050; // @[AxiLoadQueue.scala 329:31:@42155.4]
  assign loadCompleting_6 = _T_98051 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42156.4]
  assign _T_98062 = outputPriorityPorts_0_7 & dataKnown_7; // @[AxiLoadQueue.scala 328:108:@42161.4]
  assign _T_98064 = loadCompleted_7 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42162.4]
  assign _T_98065 = _T_98062 & _T_98064; // @[AxiLoadQueue.scala 329:31:@42163.4]
  assign loadCompleting_7 = _T_98065 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42164.4]
  assign _T_98076 = outputPriorityPorts_0_8 & dataKnown_8; // @[AxiLoadQueue.scala 328:108:@42169.4]
  assign _T_98078 = loadCompleted_8 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42170.4]
  assign _T_98079 = _T_98076 & _T_98078; // @[AxiLoadQueue.scala 329:31:@42171.4]
  assign loadCompleting_8 = _T_98079 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42172.4]
  assign _T_98090 = outputPriorityPorts_0_9 & dataKnown_9; // @[AxiLoadQueue.scala 328:108:@42177.4]
  assign _T_98092 = loadCompleted_9 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42178.4]
  assign _T_98093 = _T_98090 & _T_98092; // @[AxiLoadQueue.scala 329:31:@42179.4]
  assign loadCompleting_9 = _T_98093 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42180.4]
  assign _T_98104 = outputPriorityPorts_0_10 & dataKnown_10; // @[AxiLoadQueue.scala 328:108:@42185.4]
  assign _T_98106 = loadCompleted_10 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42186.4]
  assign _T_98107 = _T_98104 & _T_98106; // @[AxiLoadQueue.scala 329:31:@42187.4]
  assign loadCompleting_10 = _T_98107 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42188.4]
  assign _T_98118 = outputPriorityPorts_0_11 & dataKnown_11; // @[AxiLoadQueue.scala 328:108:@42193.4]
  assign _T_98120 = loadCompleted_11 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42194.4]
  assign _T_98121 = _T_98118 & _T_98120; // @[AxiLoadQueue.scala 329:31:@42195.4]
  assign loadCompleting_11 = _T_98121 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42196.4]
  assign _T_98132 = outputPriorityPorts_0_12 & dataKnown_12; // @[AxiLoadQueue.scala 328:108:@42201.4]
  assign _T_98134 = loadCompleted_12 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42202.4]
  assign _T_98135 = _T_98132 & _T_98134; // @[AxiLoadQueue.scala 329:31:@42203.4]
  assign loadCompleting_12 = _T_98135 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42204.4]
  assign _T_98146 = outputPriorityPorts_0_13 & dataKnown_13; // @[AxiLoadQueue.scala 328:108:@42209.4]
  assign _T_98148 = loadCompleted_13 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42210.4]
  assign _T_98149 = _T_98146 & _T_98148; // @[AxiLoadQueue.scala 329:31:@42211.4]
  assign loadCompleting_13 = _T_98149 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42212.4]
  assign _T_98160 = outputPriorityPorts_0_14 & dataKnown_14; // @[AxiLoadQueue.scala 328:108:@42217.4]
  assign _T_98162 = loadCompleted_14 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42218.4]
  assign _T_98163 = _T_98160 & _T_98162; // @[AxiLoadQueue.scala 329:31:@42219.4]
  assign loadCompleting_14 = _T_98163 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42220.4]
  assign _T_98174 = outputPriorityPorts_0_15 & dataKnown_15; // @[AxiLoadQueue.scala 328:108:@42225.4]
  assign _T_98176 = loadCompleted_15 == 1'h0; // @[AxiLoadQueue.scala 329:34:@42226.4]
  assign _T_98177 = _T_98174 & _T_98176; // @[AxiLoadQueue.scala 329:31:@42227.4]
  assign loadCompleting_15 = _T_98177 & io_loadPorts_0_ready; // @[AxiLoadQueue.scala 329:63:@42228.4]
  assign _GEN_2192 = loadCompleting_0 ? 1'h1 : loadCompleted_0; // @[AxiLoadQueue.scala 339:46:@42237.6]
  assign _GEN_2193 = initBits_0 ? 1'h0 : _GEN_2192; // @[AxiLoadQueue.scala 337:34:@42233.4]
  assign _GEN_2194 = loadCompleting_1 ? 1'h1 : loadCompleted_1; // @[AxiLoadQueue.scala 339:46:@42244.6]
  assign _GEN_2195 = initBits_1 ? 1'h0 : _GEN_2194; // @[AxiLoadQueue.scala 337:34:@42240.4]
  assign _GEN_2196 = loadCompleting_2 ? 1'h1 : loadCompleted_2; // @[AxiLoadQueue.scala 339:46:@42251.6]
  assign _GEN_2197 = initBits_2 ? 1'h0 : _GEN_2196; // @[AxiLoadQueue.scala 337:34:@42247.4]
  assign _GEN_2198 = loadCompleting_3 ? 1'h1 : loadCompleted_3; // @[AxiLoadQueue.scala 339:46:@42258.6]
  assign _GEN_2199 = initBits_3 ? 1'h0 : _GEN_2198; // @[AxiLoadQueue.scala 337:34:@42254.4]
  assign _GEN_2200 = loadCompleting_4 ? 1'h1 : loadCompleted_4; // @[AxiLoadQueue.scala 339:46:@42265.6]
  assign _GEN_2201 = initBits_4 ? 1'h0 : _GEN_2200; // @[AxiLoadQueue.scala 337:34:@42261.4]
  assign _GEN_2202 = loadCompleting_5 ? 1'h1 : loadCompleted_5; // @[AxiLoadQueue.scala 339:46:@42272.6]
  assign _GEN_2203 = initBits_5 ? 1'h0 : _GEN_2202; // @[AxiLoadQueue.scala 337:34:@42268.4]
  assign _GEN_2204 = loadCompleting_6 ? 1'h1 : loadCompleted_6; // @[AxiLoadQueue.scala 339:46:@42279.6]
  assign _GEN_2205 = initBits_6 ? 1'h0 : _GEN_2204; // @[AxiLoadQueue.scala 337:34:@42275.4]
  assign _GEN_2206 = loadCompleting_7 ? 1'h1 : loadCompleted_7; // @[AxiLoadQueue.scala 339:46:@42286.6]
  assign _GEN_2207 = initBits_7 ? 1'h0 : _GEN_2206; // @[AxiLoadQueue.scala 337:34:@42282.4]
  assign _GEN_2208 = loadCompleting_8 ? 1'h1 : loadCompleted_8; // @[AxiLoadQueue.scala 339:46:@42293.6]
  assign _GEN_2209 = initBits_8 ? 1'h0 : _GEN_2208; // @[AxiLoadQueue.scala 337:34:@42289.4]
  assign _GEN_2210 = loadCompleting_9 ? 1'h1 : loadCompleted_9; // @[AxiLoadQueue.scala 339:46:@42300.6]
  assign _GEN_2211 = initBits_9 ? 1'h0 : _GEN_2210; // @[AxiLoadQueue.scala 337:34:@42296.4]
  assign _GEN_2212 = loadCompleting_10 ? 1'h1 : loadCompleted_10; // @[AxiLoadQueue.scala 339:46:@42307.6]
  assign _GEN_2213 = initBits_10 ? 1'h0 : _GEN_2212; // @[AxiLoadQueue.scala 337:34:@42303.4]
  assign _GEN_2214 = loadCompleting_11 ? 1'h1 : loadCompleted_11; // @[AxiLoadQueue.scala 339:46:@42314.6]
  assign _GEN_2215 = initBits_11 ? 1'h0 : _GEN_2214; // @[AxiLoadQueue.scala 337:34:@42310.4]
  assign _GEN_2216 = loadCompleting_12 ? 1'h1 : loadCompleted_12; // @[AxiLoadQueue.scala 339:46:@42321.6]
  assign _GEN_2217 = initBits_12 ? 1'h0 : _GEN_2216; // @[AxiLoadQueue.scala 337:34:@42317.4]
  assign _GEN_2218 = loadCompleting_13 ? 1'h1 : loadCompleted_13; // @[AxiLoadQueue.scala 339:46:@42328.6]
  assign _GEN_2219 = initBits_13 ? 1'h0 : _GEN_2218; // @[AxiLoadQueue.scala 337:34:@42324.4]
  assign _GEN_2220 = loadCompleting_14 ? 1'h1 : loadCompleted_14; // @[AxiLoadQueue.scala 339:46:@42335.6]
  assign _GEN_2221 = initBits_14 ? 1'h0 : _GEN_2220; // @[AxiLoadQueue.scala 337:34:@42331.4]
  assign _GEN_2222 = loadCompleting_15 ? 1'h1 : loadCompleted_15; // @[AxiLoadQueue.scala 339:46:@42342.6]
  assign _GEN_2223 = initBits_15 ? 1'h0 : _GEN_2222; // @[AxiLoadQueue.scala 337:34:@42338.4]
  assign _T_98308 = _T_97967 | _T_97981; // @[AxiLoadQueue.scala 350:24:@42411.4]
  assign _T_98309 = _T_98308 | _T_97995; // @[AxiLoadQueue.scala 350:24:@42412.4]
  assign _T_98310 = _T_98309 | _T_98009; // @[AxiLoadQueue.scala 350:24:@42413.4]
  assign _T_98311 = _T_98310 | _T_98023; // @[AxiLoadQueue.scala 350:24:@42414.4]
  assign _T_98312 = _T_98311 | _T_98037; // @[AxiLoadQueue.scala 350:24:@42415.4]
  assign _T_98313 = _T_98312 | _T_98051; // @[AxiLoadQueue.scala 350:24:@42416.4]
  assign _T_98314 = _T_98313 | _T_98065; // @[AxiLoadQueue.scala 350:24:@42417.4]
  assign _T_98315 = _T_98314 | _T_98079; // @[AxiLoadQueue.scala 350:24:@42418.4]
  assign _T_98316 = _T_98315 | _T_98093; // @[AxiLoadQueue.scala 350:24:@42419.4]
  assign _T_98317 = _T_98316 | _T_98107; // @[AxiLoadQueue.scala 350:24:@42420.4]
  assign _T_98318 = _T_98317 | _T_98121; // @[AxiLoadQueue.scala 350:24:@42421.4]
  assign _T_98319 = _T_98318 | _T_98135; // @[AxiLoadQueue.scala 350:24:@42422.4]
  assign _T_98320 = _T_98319 | _T_98149; // @[AxiLoadQueue.scala 350:24:@42423.4]
  assign _T_98321 = _T_98320 | _T_98163; // @[AxiLoadQueue.scala 350:24:@42424.4]
  assign _T_98322 = _T_98321 | _T_98177; // @[AxiLoadQueue.scala 350:24:@42425.4]
  assign _T_98339 = _T_98163 ? 4'he : 4'hf; // @[Mux.scala 31:69:@42427.6]
  assign _T_98340 = _T_98149 ? 4'hd : _T_98339; // @[Mux.scala 31:69:@42428.6]
  assign _T_98341 = _T_98135 ? 4'hc : _T_98340; // @[Mux.scala 31:69:@42429.6]
  assign _T_98342 = _T_98121 ? 4'hb : _T_98341; // @[Mux.scala 31:69:@42430.6]
  assign _T_98343 = _T_98107 ? 4'ha : _T_98342; // @[Mux.scala 31:69:@42431.6]
  assign _T_98344 = _T_98093 ? 4'h9 : _T_98343; // @[Mux.scala 31:69:@42432.6]
  assign _T_98345 = _T_98079 ? 4'h8 : _T_98344; // @[Mux.scala 31:69:@42433.6]
  assign _T_98346 = _T_98065 ? 4'h7 : _T_98345; // @[Mux.scala 31:69:@42434.6]
  assign _T_98347 = _T_98051 ? 4'h6 : _T_98346; // @[Mux.scala 31:69:@42435.6]
  assign _T_98348 = _T_98037 ? 4'h5 : _T_98347; // @[Mux.scala 31:69:@42436.6]
  assign _T_98349 = _T_98023 ? 4'h4 : _T_98348; // @[Mux.scala 31:69:@42437.6]
  assign _T_98350 = _T_98009 ? 4'h3 : _T_98349; // @[Mux.scala 31:69:@42438.6]
  assign _T_98351 = _T_97995 ? 4'h2 : _T_98350; // @[Mux.scala 31:69:@42439.6]
  assign _T_98352 = _T_97981 ? 4'h1 : _T_98351; // @[Mux.scala 31:69:@42440.6]
  assign _T_98353 = _T_97967 ? 4'h0 : _T_98352; // @[Mux.scala 31:69:@42441.6]
  assign _GEN_2225 = 4'h1 == _T_98353 ? dataQ_1 : dataQ_0; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2226 = 4'h2 == _T_98353 ? dataQ_2 : _GEN_2225; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2227 = 4'h3 == _T_98353 ? dataQ_3 : _GEN_2226; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2228 = 4'h4 == _T_98353 ? dataQ_4 : _GEN_2227; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2229 = 4'h5 == _T_98353 ? dataQ_5 : _GEN_2228; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2230 = 4'h6 == _T_98353 ? dataQ_6 : _GEN_2229; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2231 = 4'h7 == _T_98353 ? dataQ_7 : _GEN_2230; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2232 = 4'h8 == _T_98353 ? dataQ_8 : _GEN_2231; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2233 = 4'h9 == _T_98353 ? dataQ_9 : _GEN_2232; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2234 = 4'ha == _T_98353 ? dataQ_10 : _GEN_2233; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2235 = 4'hb == _T_98353 ? dataQ_11 : _GEN_2234; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2236 = 4'hc == _T_98353 ? dataQ_12 : _GEN_2235; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2237 = 4'hd == _T_98353 ? dataQ_13 : _GEN_2236; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2238 = 4'he == _T_98353 ? dataQ_14 : _GEN_2237; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2239 = 4'hf == _T_98353 ? dataQ_15 : _GEN_2238; // @[AxiLoadQueue.scala 351:37:@42442.6]
  assign _GEN_2243 = 4'h1 == head ? loadCompleted_1 : loadCompleted_0; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2244 = 4'h2 == head ? loadCompleted_2 : _GEN_2243; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2245 = 4'h3 == head ? loadCompleted_3 : _GEN_2244; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2246 = 4'h4 == head ? loadCompleted_4 : _GEN_2245; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2247 = 4'h5 == head ? loadCompleted_5 : _GEN_2246; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2248 = 4'h6 == head ? loadCompleted_6 : _GEN_2247; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2249 = 4'h7 == head ? loadCompleted_7 : _GEN_2248; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2250 = 4'h8 == head ? loadCompleted_8 : _GEN_2249; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2251 = 4'h9 == head ? loadCompleted_9 : _GEN_2250; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2252 = 4'ha == head ? loadCompleted_10 : _GEN_2251; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2253 = 4'hb == head ? loadCompleted_11 : _GEN_2252; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2254 = 4'hc == head ? loadCompleted_12 : _GEN_2253; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2255 = 4'hd == head ? loadCompleted_13 : _GEN_2254; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2256 = 4'he == head ? loadCompleted_14 : _GEN_2255; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2257 = 4'hf == head ? loadCompleted_15 : _GEN_2256; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2259 = 4'h1 == head ? loadCompleting_1 : loadCompleting_0; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2260 = 4'h2 == head ? loadCompleting_2 : _GEN_2259; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2261 = 4'h3 == head ? loadCompleting_3 : _GEN_2260; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2262 = 4'h4 == head ? loadCompleting_4 : _GEN_2261; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2263 = 4'h5 == head ? loadCompleting_5 : _GEN_2262; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2264 = 4'h6 == head ? loadCompleting_6 : _GEN_2263; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2265 = 4'h7 == head ? loadCompleting_7 : _GEN_2264; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2266 = 4'h8 == head ? loadCompleting_8 : _GEN_2265; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2267 = 4'h9 == head ? loadCompleting_9 : _GEN_2266; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2268 = 4'ha == head ? loadCompleting_10 : _GEN_2267; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2269 = 4'hb == head ? loadCompleting_11 : _GEN_2268; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2270 = 4'hc == head ? loadCompleting_12 : _GEN_2269; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2271 = 4'hd == head ? loadCompleting_13 : _GEN_2270; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2272 = 4'he == head ? loadCompleting_14 : _GEN_2271; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _GEN_2273 = 4'hf == head ? loadCompleting_15 : _GEN_2272; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _T_98364 = _GEN_2257 | _GEN_2273; // @[AxiLoadQueue.scala 365:29:@42449.4]
  assign _T_98365 = head != tail; // @[AxiLoadQueue.scala 365:63:@42450.4]
  assign _T_98367 = io_loadEmpty == 1'h0; // @[AxiLoadQueue.scala 365:75:@42451.4]
  assign _T_98368 = _T_98365 | _T_98367; // @[AxiLoadQueue.scala 365:72:@42452.4]
  assign _T_98369 = _T_98364 & _T_98368; // @[AxiLoadQueue.scala 365:54:@42453.4]
  assign _T_98372 = head + 4'h1; // @[util.scala 10:8:@42455.6]
  assign _GEN_64 = _T_98372 % 5'h10; // @[util.scala 10:14:@42456.6]
  assign _T_98373 = _GEN_64[4:0]; // @[util.scala 10:14:@42456.6]
  assign _GEN_2274 = _T_98369 ? _T_98373 : {{1'd0}, head}; // @[AxiLoadQueue.scala 365:91:@42454.4]
  assign _GEN_2372 = {{3'd0}, io_bbNumLoads}; // @[util.scala 10:8:@42460.6]
  assign _T_98375 = tail + _GEN_2372; // @[util.scala 10:8:@42460.6]
  assign _GEN_65 = _T_98375 % 5'h10; // @[util.scala 10:14:@42461.6]
  assign _T_98376 = _GEN_65[4:0]; // @[util.scala 10:14:@42461.6]
  assign _GEN_2275 = io_bbStart ? _T_98376 : {{1'd0}, tail}; // @[AxiLoadQueue.scala 369:20:@42459.4]
  assign _T_98378 = allocatedEntries_0 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42464.4]
  assign _T_98379 = loadCompleted_0 | _T_98378; // @[AxiLoadQueue.scala 373:79:@42465.4]
  assign _T_98381 = allocatedEntries_1 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42466.4]
  assign _T_98382 = loadCompleted_1 | _T_98381; // @[AxiLoadQueue.scala 373:79:@42467.4]
  assign _T_98384 = allocatedEntries_2 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42468.4]
  assign _T_98385 = loadCompleted_2 | _T_98384; // @[AxiLoadQueue.scala 373:79:@42469.4]
  assign _T_98387 = allocatedEntries_3 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42470.4]
  assign _T_98388 = loadCompleted_3 | _T_98387; // @[AxiLoadQueue.scala 373:79:@42471.4]
  assign _T_98390 = allocatedEntries_4 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42472.4]
  assign _T_98391 = loadCompleted_4 | _T_98390; // @[AxiLoadQueue.scala 373:79:@42473.4]
  assign _T_98393 = allocatedEntries_5 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42474.4]
  assign _T_98394 = loadCompleted_5 | _T_98393; // @[AxiLoadQueue.scala 373:79:@42475.4]
  assign _T_98396 = allocatedEntries_6 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42476.4]
  assign _T_98397 = loadCompleted_6 | _T_98396; // @[AxiLoadQueue.scala 373:79:@42477.4]
  assign _T_98399 = allocatedEntries_7 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42478.4]
  assign _T_98400 = loadCompleted_7 | _T_98399; // @[AxiLoadQueue.scala 373:79:@42479.4]
  assign _T_98402 = allocatedEntries_8 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42480.4]
  assign _T_98403 = loadCompleted_8 | _T_98402; // @[AxiLoadQueue.scala 373:79:@42481.4]
  assign _T_98405 = allocatedEntries_9 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42482.4]
  assign _T_98406 = loadCompleted_9 | _T_98405; // @[AxiLoadQueue.scala 373:79:@42483.4]
  assign _T_98408 = allocatedEntries_10 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42484.4]
  assign _T_98409 = loadCompleted_10 | _T_98408; // @[AxiLoadQueue.scala 373:79:@42485.4]
  assign _T_98411 = allocatedEntries_11 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42486.4]
  assign _T_98412 = loadCompleted_11 | _T_98411; // @[AxiLoadQueue.scala 373:79:@42487.4]
  assign _T_98414 = allocatedEntries_12 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42488.4]
  assign _T_98415 = loadCompleted_12 | _T_98414; // @[AxiLoadQueue.scala 373:79:@42489.4]
  assign _T_98417 = allocatedEntries_13 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42490.4]
  assign _T_98418 = loadCompleted_13 | _T_98417; // @[AxiLoadQueue.scala 373:79:@42491.4]
  assign _T_98420 = allocatedEntries_14 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42492.4]
  assign _T_98421 = loadCompleted_14 | _T_98420; // @[AxiLoadQueue.scala 373:79:@42493.4]
  assign _T_98423 = allocatedEntries_15 == 1'h0; // @[AxiLoadQueue.scala 373:82:@42494.4]
  assign _T_98424 = loadCompleted_15 | _T_98423; // @[AxiLoadQueue.scala 373:79:@42495.4]
  assign _T_98449 = _T_98379 & _T_98382; // @[AxiLoadQueue.scala 373:96:@42514.4]
  assign _T_98450 = _T_98449 & _T_98385; // @[AxiLoadQueue.scala 373:96:@42515.4]
  assign _T_98451 = _T_98450 & _T_98388; // @[AxiLoadQueue.scala 373:96:@42516.4]
  assign _T_98452 = _T_98451 & _T_98391; // @[AxiLoadQueue.scala 373:96:@42517.4]
  assign _T_98453 = _T_98452 & _T_98394; // @[AxiLoadQueue.scala 373:96:@42518.4]
  assign _T_98454 = _T_98453 & _T_98397; // @[AxiLoadQueue.scala 373:96:@42519.4]
  assign _T_98455 = _T_98454 & _T_98400; // @[AxiLoadQueue.scala 373:96:@42520.4]
  assign _T_98456 = _T_98455 & _T_98403; // @[AxiLoadQueue.scala 373:96:@42521.4]
  assign _T_98457 = _T_98456 & _T_98406; // @[AxiLoadQueue.scala 373:96:@42522.4]
  assign _T_98458 = _T_98457 & _T_98409; // @[AxiLoadQueue.scala 373:96:@42523.4]
  assign _T_98459 = _T_98458 & _T_98412; // @[AxiLoadQueue.scala 373:96:@42524.4]
  assign _T_98460 = _T_98459 & _T_98415; // @[AxiLoadQueue.scala 373:96:@42525.4]
  assign _T_98461 = _T_98460 & _T_98418; // @[AxiLoadQueue.scala 373:96:@42526.4]
  assign _T_98462 = _T_98461 & _T_98421; // @[AxiLoadQueue.scala 373:96:@42527.4]
  assign io_loadTail = tail; // @[AxiLoadQueue.scala 382:15:@42531.4]
  assign io_loadHead = head; // @[AxiLoadQueue.scala 381:15:@42530.4]
  assign io_loadEmpty = _T_98462 & _T_98424; // @[AxiLoadQueue.scala 373:16:@42529.4]
  assign io_loadAddrDone_0 = addrKnown_0; // @[AxiLoadQueue.scala 384:19:@42548.4]
  assign io_loadAddrDone_1 = addrKnown_1; // @[AxiLoadQueue.scala 384:19:@42549.4]
  assign io_loadAddrDone_2 = addrKnown_2; // @[AxiLoadQueue.scala 384:19:@42550.4]
  assign io_loadAddrDone_3 = addrKnown_3; // @[AxiLoadQueue.scala 384:19:@42551.4]
  assign io_loadAddrDone_4 = addrKnown_4; // @[AxiLoadQueue.scala 384:19:@42552.4]
  assign io_loadAddrDone_5 = addrKnown_5; // @[AxiLoadQueue.scala 384:19:@42553.4]
  assign io_loadAddrDone_6 = addrKnown_6; // @[AxiLoadQueue.scala 384:19:@42554.4]
  assign io_loadAddrDone_7 = addrKnown_7; // @[AxiLoadQueue.scala 384:19:@42555.4]
  assign io_loadAddrDone_8 = addrKnown_8; // @[AxiLoadQueue.scala 384:19:@42556.4]
  assign io_loadAddrDone_9 = addrKnown_9; // @[AxiLoadQueue.scala 384:19:@42557.4]
  assign io_loadAddrDone_10 = addrKnown_10; // @[AxiLoadQueue.scala 384:19:@42558.4]
  assign io_loadAddrDone_11 = addrKnown_11; // @[AxiLoadQueue.scala 384:19:@42559.4]
  assign io_loadAddrDone_12 = addrKnown_12; // @[AxiLoadQueue.scala 384:19:@42560.4]
  assign io_loadAddrDone_13 = addrKnown_13; // @[AxiLoadQueue.scala 384:19:@42561.4]
  assign io_loadAddrDone_14 = addrKnown_14; // @[AxiLoadQueue.scala 384:19:@42562.4]
  assign io_loadAddrDone_15 = addrKnown_15; // @[AxiLoadQueue.scala 384:19:@42563.4]
  assign io_loadDataDone_0 = dataKnown_0; // @[AxiLoadQueue.scala 385:19:@42564.4]
  assign io_loadDataDone_1 = dataKnown_1; // @[AxiLoadQueue.scala 385:19:@42565.4]
  assign io_loadDataDone_2 = dataKnown_2; // @[AxiLoadQueue.scala 385:19:@42566.4]
  assign io_loadDataDone_3 = dataKnown_3; // @[AxiLoadQueue.scala 385:19:@42567.4]
  assign io_loadDataDone_4 = dataKnown_4; // @[AxiLoadQueue.scala 385:19:@42568.4]
  assign io_loadDataDone_5 = dataKnown_5; // @[AxiLoadQueue.scala 385:19:@42569.4]
  assign io_loadDataDone_6 = dataKnown_6; // @[AxiLoadQueue.scala 385:19:@42570.4]
  assign io_loadDataDone_7 = dataKnown_7; // @[AxiLoadQueue.scala 385:19:@42571.4]
  assign io_loadDataDone_8 = dataKnown_8; // @[AxiLoadQueue.scala 385:19:@42572.4]
  assign io_loadDataDone_9 = dataKnown_9; // @[AxiLoadQueue.scala 385:19:@42573.4]
  assign io_loadDataDone_10 = dataKnown_10; // @[AxiLoadQueue.scala 385:19:@42574.4]
  assign io_loadDataDone_11 = dataKnown_11; // @[AxiLoadQueue.scala 385:19:@42575.4]
  assign io_loadDataDone_12 = dataKnown_12; // @[AxiLoadQueue.scala 385:19:@42576.4]
  assign io_loadDataDone_13 = dataKnown_13; // @[AxiLoadQueue.scala 385:19:@42577.4]
  assign io_loadDataDone_14 = dataKnown_14; // @[AxiLoadQueue.scala 385:19:@42578.4]
  assign io_loadDataDone_15 = dataKnown_15; // @[AxiLoadQueue.scala 385:19:@42579.4]
  assign io_loadAddrQueue_0 = addrQ_0; // @[AxiLoadQueue.scala 383:20:@42532.4]
  assign io_loadAddrQueue_1 = addrQ_1; // @[AxiLoadQueue.scala 383:20:@42533.4]
  assign io_loadAddrQueue_2 = addrQ_2; // @[AxiLoadQueue.scala 383:20:@42534.4]
  assign io_loadAddrQueue_3 = addrQ_3; // @[AxiLoadQueue.scala 383:20:@42535.4]
  assign io_loadAddrQueue_4 = addrQ_4; // @[AxiLoadQueue.scala 383:20:@42536.4]
  assign io_loadAddrQueue_5 = addrQ_5; // @[AxiLoadQueue.scala 383:20:@42537.4]
  assign io_loadAddrQueue_6 = addrQ_6; // @[AxiLoadQueue.scala 383:20:@42538.4]
  assign io_loadAddrQueue_7 = addrQ_7; // @[AxiLoadQueue.scala 383:20:@42539.4]
  assign io_loadAddrQueue_8 = addrQ_8; // @[AxiLoadQueue.scala 383:20:@42540.4]
  assign io_loadAddrQueue_9 = addrQ_9; // @[AxiLoadQueue.scala 383:20:@42541.4]
  assign io_loadAddrQueue_10 = addrQ_10; // @[AxiLoadQueue.scala 383:20:@42542.4]
  assign io_loadAddrQueue_11 = addrQ_11; // @[AxiLoadQueue.scala 383:20:@42543.4]
  assign io_loadAddrQueue_12 = addrQ_12; // @[AxiLoadQueue.scala 383:20:@42544.4]
  assign io_loadAddrQueue_13 = addrQ_13; // @[AxiLoadQueue.scala 383:20:@42545.4]
  assign io_loadAddrQueue_14 = addrQ_14; // @[AxiLoadQueue.scala 383:20:@42546.4]
  assign io_loadAddrQueue_15 = addrQ_15; // @[AxiLoadQueue.scala 383:20:@42547.4]
  assign io_loadPorts_0_valid = _T_98321 | _T_98177; // @[AxiLoadQueue.scala 352:38:@42443.6 AxiLoadQueue.scala 355:38:@42447.6]
  assign io_loadPorts_0_bits = _T_98322 ? _GEN_2239 : 32'h0; // @[AxiLoadQueue.scala 351:37:@42442.6 AxiLoadQueue.scala 354:37:@42446.6]
  assign io_loadAddrToMem = 4'hf == _T_92263 ? addrQ_15 : _GEN_1966; // @[AxiLoadQueue.scala 223:20:@37799.4]
  assign io_loadQIdxForAddrOut_valid = _T_92279 | priorityLoadRequest_15; // @[AxiLoadQueue.scala 222:31:@37783.4]
  assign io_loadQIdxForAddrOut_bits = priorityLoadRequest_0 ? 4'h0 : _T_92262; // @[AxiLoadQueue.scala 221:30:@37766.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  head = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tail = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  offsetQ_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  offsetQ_1 = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  offsetQ_2 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  offsetQ_3 = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  offsetQ_4 = _RAND_6[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  offsetQ_5 = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  offsetQ_6 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  offsetQ_7 = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  offsetQ_8 = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  offsetQ_9 = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  offsetQ_10 = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  offsetQ_11 = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  offsetQ_12 = _RAND_14[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  offsetQ_13 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  offsetQ_14 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  offsetQ_15 = _RAND_17[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  portQ_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  portQ_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  portQ_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  portQ_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  portQ_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  portQ_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  portQ_6 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  portQ_7 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  portQ_8 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  portQ_9 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  portQ_10 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  portQ_11 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  portQ_12 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  portQ_13 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  portQ_14 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  portQ_15 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  addrQ_0 = _RAND_34[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  addrQ_1 = _RAND_35[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  addrQ_2 = _RAND_36[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  addrQ_3 = _RAND_37[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  addrQ_4 = _RAND_38[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  addrQ_5 = _RAND_39[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  addrQ_6 = _RAND_40[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  addrQ_7 = _RAND_41[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  addrQ_8 = _RAND_42[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  addrQ_9 = _RAND_43[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  addrQ_10 = _RAND_44[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  addrQ_11 = _RAND_45[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  addrQ_12 = _RAND_46[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  addrQ_13 = _RAND_47[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  addrQ_14 = _RAND_48[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  addrQ_15 = _RAND_49[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  dataQ_0 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  dataQ_1 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  dataQ_2 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  dataQ_3 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  dataQ_4 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  dataQ_5 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  dataQ_6 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  dataQ_7 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dataQ_8 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  dataQ_9 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  dataQ_10 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  dataQ_11 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  dataQ_12 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  dataQ_13 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  dataQ_14 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  dataQ_15 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  addrKnown_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  addrKnown_1 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  addrKnown_2 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  addrKnown_3 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  addrKnown_4 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  addrKnown_5 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  addrKnown_6 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  addrKnown_7 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  addrKnown_8 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  addrKnown_9 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  addrKnown_10 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  addrKnown_11 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  addrKnown_12 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  addrKnown_13 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  addrKnown_14 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  addrKnown_15 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataKnown_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  dataKnown_1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  dataKnown_2 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  dataKnown_3 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  dataKnown_4 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dataKnown_5 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dataKnown_6 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dataKnown_7 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dataKnown_8 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dataKnown_9 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dataKnown_10 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dataKnown_11 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dataKnown_12 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dataKnown_13 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dataKnown_14 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dataKnown_15 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  loadCompleted_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  loadCompleted_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  loadCompleted_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  loadCompleted_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  loadCompleted_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  loadCompleted_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  loadCompleted_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  loadCompleted_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  loadCompleted_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  loadCompleted_9 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  loadCompleted_10 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  loadCompleted_11 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  loadCompleted_12 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  loadCompleted_13 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  loadCompleted_14 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  loadCompleted_15 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  allocatedEntries_0 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  allocatedEntries_1 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  allocatedEntries_2 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  allocatedEntries_3 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  allocatedEntries_4 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  allocatedEntries_5 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  allocatedEntries_6 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  allocatedEntries_7 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  allocatedEntries_8 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  allocatedEntries_9 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  allocatedEntries_10 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  allocatedEntries_11 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  allocatedEntries_12 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  allocatedEntries_13 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  allocatedEntries_14 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  allocatedEntries_15 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  bypassInitiated_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  bypassInitiated_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  bypassInitiated_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  bypassInitiated_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  bypassInitiated_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  bypassInitiated_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  bypassInitiated_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  bypassInitiated_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  bypassInitiated_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  bypassInitiated_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  bypassInitiated_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  bypassInitiated_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  bypassInitiated_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  bypassInitiated_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  bypassInitiated_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  bypassInitiated_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  checkBits_0 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  checkBits_1 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  checkBits_2 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  checkBits_3 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  checkBits_4 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  checkBits_5 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  checkBits_6 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  checkBits_7 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  checkBits_8 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  checkBits_9 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  checkBits_10 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  checkBits_11 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  checkBits_12 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  checkBits_13 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  checkBits_14 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  checkBits_15 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  previousStoreHead = _RAND_162[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  conflictPReg_0_0 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  conflictPReg_0_1 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  conflictPReg_0_2 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  conflictPReg_0_3 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  conflictPReg_0_4 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  conflictPReg_0_5 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  conflictPReg_0_6 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  conflictPReg_0_7 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  conflictPReg_0_8 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  conflictPReg_0_9 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  conflictPReg_0_10 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  conflictPReg_0_11 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  conflictPReg_0_12 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  conflictPReg_0_13 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  conflictPReg_0_14 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  conflictPReg_0_15 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  conflictPReg_1_0 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  conflictPReg_1_1 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  conflictPReg_1_2 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  conflictPReg_1_3 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  conflictPReg_1_4 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  conflictPReg_1_5 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  conflictPReg_1_6 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  conflictPReg_1_7 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  conflictPReg_1_8 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  conflictPReg_1_9 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  conflictPReg_1_10 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  conflictPReg_1_11 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  conflictPReg_1_12 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  conflictPReg_1_13 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  conflictPReg_1_14 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  conflictPReg_1_15 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  conflictPReg_2_0 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  conflictPReg_2_1 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  conflictPReg_2_2 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  conflictPReg_2_3 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  conflictPReg_2_4 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  conflictPReg_2_5 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  conflictPReg_2_6 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  conflictPReg_2_7 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  conflictPReg_2_8 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  conflictPReg_2_9 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  conflictPReg_2_10 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  conflictPReg_2_11 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  conflictPReg_2_12 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  conflictPReg_2_13 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  conflictPReg_2_14 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  conflictPReg_2_15 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  conflictPReg_3_0 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  conflictPReg_3_1 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  conflictPReg_3_2 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  conflictPReg_3_3 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  conflictPReg_3_4 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  conflictPReg_3_5 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  conflictPReg_3_6 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  conflictPReg_3_7 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  conflictPReg_3_8 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  conflictPReg_3_9 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  conflictPReg_3_10 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  conflictPReg_3_11 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  conflictPReg_3_12 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  conflictPReg_3_13 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  conflictPReg_3_14 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  conflictPReg_3_15 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  conflictPReg_4_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  conflictPReg_4_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  conflictPReg_4_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  conflictPReg_4_3 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  conflictPReg_4_4 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  conflictPReg_4_5 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  conflictPReg_4_6 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  conflictPReg_4_7 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  conflictPReg_4_8 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  conflictPReg_4_9 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  conflictPReg_4_10 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  conflictPReg_4_11 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  conflictPReg_4_12 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  conflictPReg_4_13 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  conflictPReg_4_14 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  conflictPReg_4_15 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  conflictPReg_5_0 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  conflictPReg_5_1 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  conflictPReg_5_2 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  conflictPReg_5_3 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  conflictPReg_5_4 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  conflictPReg_5_5 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  conflictPReg_5_6 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  conflictPReg_5_7 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  conflictPReg_5_8 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  conflictPReg_5_9 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  conflictPReg_5_10 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  conflictPReg_5_11 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  conflictPReg_5_12 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  conflictPReg_5_13 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  conflictPReg_5_14 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  conflictPReg_5_15 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  conflictPReg_6_0 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  conflictPReg_6_1 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  conflictPReg_6_2 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  conflictPReg_6_3 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  conflictPReg_6_4 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  conflictPReg_6_5 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  conflictPReg_6_6 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  conflictPReg_6_7 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  conflictPReg_6_8 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  conflictPReg_6_9 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  conflictPReg_6_10 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  conflictPReg_6_11 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  conflictPReg_6_12 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  conflictPReg_6_13 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  conflictPReg_6_14 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  conflictPReg_6_15 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  conflictPReg_7_0 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  conflictPReg_7_1 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  conflictPReg_7_2 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  conflictPReg_7_3 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  conflictPReg_7_4 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  conflictPReg_7_5 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  conflictPReg_7_6 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  conflictPReg_7_7 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  conflictPReg_7_8 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  conflictPReg_7_9 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  conflictPReg_7_10 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  conflictPReg_7_11 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  conflictPReg_7_12 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  conflictPReg_7_13 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  conflictPReg_7_14 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  conflictPReg_7_15 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  conflictPReg_8_0 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  conflictPReg_8_1 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  conflictPReg_8_2 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  conflictPReg_8_3 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  conflictPReg_8_4 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  conflictPReg_8_5 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  conflictPReg_8_6 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  conflictPReg_8_7 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  conflictPReg_8_8 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  conflictPReg_8_9 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  conflictPReg_8_10 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  conflictPReg_8_11 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  conflictPReg_8_12 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  conflictPReg_8_13 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  conflictPReg_8_14 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  conflictPReg_8_15 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  conflictPReg_9_0 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  conflictPReg_9_1 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  conflictPReg_9_2 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  conflictPReg_9_3 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  conflictPReg_9_4 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  conflictPReg_9_5 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  conflictPReg_9_6 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  conflictPReg_9_7 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  conflictPReg_9_8 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  conflictPReg_9_9 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  conflictPReg_9_10 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  conflictPReg_9_11 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  conflictPReg_9_12 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  conflictPReg_9_13 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  conflictPReg_9_14 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  conflictPReg_9_15 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  conflictPReg_10_0 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  conflictPReg_10_1 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  conflictPReg_10_2 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  conflictPReg_10_3 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  conflictPReg_10_4 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  conflictPReg_10_5 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  conflictPReg_10_6 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  conflictPReg_10_7 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  conflictPReg_10_8 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  conflictPReg_10_9 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  conflictPReg_10_10 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  conflictPReg_10_11 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  conflictPReg_10_12 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  conflictPReg_10_13 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  conflictPReg_10_14 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  conflictPReg_10_15 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  conflictPReg_11_0 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  conflictPReg_11_1 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  conflictPReg_11_2 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  conflictPReg_11_3 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  conflictPReg_11_4 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  conflictPReg_11_5 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  conflictPReg_11_6 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  conflictPReg_11_7 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  conflictPReg_11_8 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  conflictPReg_11_9 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  conflictPReg_11_10 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  conflictPReg_11_11 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  conflictPReg_11_12 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  conflictPReg_11_13 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  conflictPReg_11_14 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  conflictPReg_11_15 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  conflictPReg_12_0 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  conflictPReg_12_1 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  conflictPReg_12_2 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  conflictPReg_12_3 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  conflictPReg_12_4 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  conflictPReg_12_5 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  conflictPReg_12_6 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  conflictPReg_12_7 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  conflictPReg_12_8 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  conflictPReg_12_9 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  conflictPReg_12_10 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  conflictPReg_12_11 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  conflictPReg_12_12 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  conflictPReg_12_13 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  conflictPReg_12_14 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  conflictPReg_12_15 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  conflictPReg_13_0 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  conflictPReg_13_1 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  conflictPReg_13_2 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  conflictPReg_13_3 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  conflictPReg_13_4 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  conflictPReg_13_5 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  conflictPReg_13_6 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  conflictPReg_13_7 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  conflictPReg_13_8 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  conflictPReg_13_9 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  conflictPReg_13_10 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  conflictPReg_13_11 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  conflictPReg_13_12 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  conflictPReg_13_13 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  conflictPReg_13_14 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  conflictPReg_13_15 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  conflictPReg_14_0 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  conflictPReg_14_1 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  conflictPReg_14_2 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  conflictPReg_14_3 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  conflictPReg_14_4 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  conflictPReg_14_5 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  conflictPReg_14_6 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  conflictPReg_14_7 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  conflictPReg_14_8 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  conflictPReg_14_9 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  conflictPReg_14_10 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  conflictPReg_14_11 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  conflictPReg_14_12 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  conflictPReg_14_13 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  conflictPReg_14_14 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  conflictPReg_14_15 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  conflictPReg_15_0 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  conflictPReg_15_1 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  conflictPReg_15_2 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  conflictPReg_15_3 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  conflictPReg_15_4 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  conflictPReg_15_5 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  conflictPReg_15_6 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  conflictPReg_15_7 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  conflictPReg_15_8 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  conflictPReg_15_9 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  conflictPReg_15_10 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  conflictPReg_15_11 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  conflictPReg_15_12 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  conflictPReg_15_13 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  conflictPReg_15_14 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  conflictPReg_15_15 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_0 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_1 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_2 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_3 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_4 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_5 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_6 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_7 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_8 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_9 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_10 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_11 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_12 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_13 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_14 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_0_15 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_0 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_1 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_2 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_3 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_4 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_5 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_6 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_7 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_8 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_9 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_10 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_11 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_12 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_13 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_14 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_1_15 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_0 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_1 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_2 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_3 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_4 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_5 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_6 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_7 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_8 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_9 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_10 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_11 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_12 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_13 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_14 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_2_15 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_0 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_1 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_2 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_3 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_4 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_5 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_6 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_7 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_8 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_9 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_10 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_11 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_12 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_13 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_14 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_3_15 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_0 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_1 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_2 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_3 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_4 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_5 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_6 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_7 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_8 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_9 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_10 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_11 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_12 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_13 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_14 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_4_15 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_0 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_1 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_2 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_3 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_4 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_5 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_6 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_7 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_8 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_9 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_10 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_11 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_12 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_13 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_14 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_5_15 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_0 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_1 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_2 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_3 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_4 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_5 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_6 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_7 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_8 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_9 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_10 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_11 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_12 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_13 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_14 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_6_15 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_0 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_1 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_2 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_3 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_4 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_5 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_6 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_7 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_8 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_9 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_10 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_11 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_12 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_13 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_14 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_7_15 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_0 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_1 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_2 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_3 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_4 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_5 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_6 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_7 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_8 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_9 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_10 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_11 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_12 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_13 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_14 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_8_15 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_0 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_1 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_2 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_3 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_4 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_5 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_6 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_7 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_8 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_9 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_10 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_11 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_12 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_13 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_14 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_9_15 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_0 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_1 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_2 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_3 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_4 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_5 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_6 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_7 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_8 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_9 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_10 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_11 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_12 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_13 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_14 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_10_15 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_0 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_1 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_2 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_3 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_4 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_5 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_6 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_7 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_8 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_9 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_10 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_11 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_12 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_13 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_14 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_11_15 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_0 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_1 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_2 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_3 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_4 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_5 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_6 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_7 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_8 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_9 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_10 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_11 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_12 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_13 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_14 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_12_15 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_0 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_1 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_2 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_3 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_4 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_5 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_6 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_7 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_8 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_9 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_10 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_11 = _RAND_638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_12 = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_13 = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_14 = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_13_15 = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_0 = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_1 = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_2 = _RAND_645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_3 = _RAND_646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_4 = _RAND_647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_5 = _RAND_648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_6 = _RAND_649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_7 = _RAND_650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_8 = _RAND_651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_9 = _RAND_652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_10 = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_11 = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_12 = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_13 = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_14 = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_14_15 = _RAND_658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_0 = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_1 = _RAND_660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_2 = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_3 = _RAND_662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_4 = _RAND_663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_5 = _RAND_664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_6 = _RAND_665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_7 = _RAND_666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_8 = _RAND_667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_9 = _RAND_668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_10 = _RAND_669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_11 = _RAND_670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_12 = _RAND_671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_13 = _RAND_672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_14 = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  storeAddrNotKnownFlagsPReg_15_15 = _RAND_674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_0 = _RAND_675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_1 = _RAND_676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_2 = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_3 = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_4 = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_5 = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_6 = _RAND_681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_7 = _RAND_682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_8 = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_9 = _RAND_684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_10 = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_11 = _RAND_686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_12 = _RAND_687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_13 = _RAND_688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_14 = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  shiftedStoreDataKnownPReg_15 = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  shiftedStoreDataQPreg_0 = _RAND_691[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  shiftedStoreDataQPreg_1 = _RAND_692[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  shiftedStoreDataQPreg_2 = _RAND_693[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  shiftedStoreDataQPreg_3 = _RAND_694[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  shiftedStoreDataQPreg_4 = _RAND_695[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  shiftedStoreDataQPreg_5 = _RAND_696[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  shiftedStoreDataQPreg_6 = _RAND_697[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  shiftedStoreDataQPreg_7 = _RAND_698[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  shiftedStoreDataQPreg_8 = _RAND_699[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  shiftedStoreDataQPreg_9 = _RAND_700[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  shiftedStoreDataQPreg_10 = _RAND_701[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  shiftedStoreDataQPreg_11 = _RAND_702[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  shiftedStoreDataQPreg_12 = _RAND_703[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  shiftedStoreDataQPreg_13 = _RAND_704[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  shiftedStoreDataQPreg_14 = _RAND_705[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  shiftedStoreDataQPreg_15 = _RAND_706[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  addrKnownPReg_0 = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  addrKnownPReg_1 = _RAND_708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  addrKnownPReg_2 = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  addrKnownPReg_3 = _RAND_710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  addrKnownPReg_4 = _RAND_711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  addrKnownPReg_5 = _RAND_712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  addrKnownPReg_6 = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  addrKnownPReg_7 = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  addrKnownPReg_8 = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  addrKnownPReg_9 = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  addrKnownPReg_10 = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  addrKnownPReg_11 = _RAND_718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  addrKnownPReg_12 = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  addrKnownPReg_13 = _RAND_720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  addrKnownPReg_14 = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  addrKnownPReg_15 = _RAND_722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  dataKnownPReg_0 = _RAND_723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  dataKnownPReg_1 = _RAND_724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  dataKnownPReg_2 = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  dataKnownPReg_3 = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  dataKnownPReg_4 = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  dataKnownPReg_5 = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  dataKnownPReg_6 = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  dataKnownPReg_7 = _RAND_730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  dataKnownPReg_8 = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  dataKnownPReg_9 = _RAND_732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  dataKnownPReg_10 = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  dataKnownPReg_11 = _RAND_734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  dataKnownPReg_12 = _RAND_735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  dataKnownPReg_13 = _RAND_736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  dataKnownPReg_14 = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  dataKnownPReg_15 = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  loadInitiated_15 = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  loadInitiated_14 = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  loadInitiated_13 = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  loadInitiated_12 = _RAND_742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  loadInitiated_11 = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  loadInitiated_10 = _RAND_744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  loadInitiated_9 = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  loadInitiated_8 = _RAND_746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  loadInitiated_7 = _RAND_747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  loadInitiated_6 = _RAND_748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  loadInitiated_5 = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  loadInitiated_4 = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  loadInitiated_3 = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  loadInitiated_2 = _RAND_752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  loadInitiated_1 = _RAND_753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  loadInitiated_0 = _RAND_754[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      head <= 4'h0;
    end else begin
      head <= _GEN_2274[3:0];
    end
    if (reset) begin
      tail <= 4'h0;
    end else begin
      tail <= _GEN_2275[3:0];
    end
    if (reset) begin
      offsetQ_0 <= 4'h0;
    end else begin
      if (initBits_0) begin
        if (4'hf == _T_1930) begin
          offsetQ_0 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1930) begin
            offsetQ_0 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1930) begin
              offsetQ_0 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1930) begin
                offsetQ_0 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1930) begin
                  offsetQ_0 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1930) begin
                    offsetQ_0 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1930) begin
                      offsetQ_0 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1930) begin
                        offsetQ_0 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1930) begin
                          offsetQ_0 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1930) begin
                            offsetQ_0 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1930) begin
                              offsetQ_0 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1930) begin
                                offsetQ_0 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1930) begin
                                  offsetQ_0 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1930) begin
                                    offsetQ_0 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1930) begin
                                      offsetQ_0 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_0 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_1 <= 4'h0;
    end else begin
      if (initBits_1) begin
        if (4'hf == _T_1948) begin
          offsetQ_1 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1948) begin
            offsetQ_1 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1948) begin
              offsetQ_1 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1948) begin
                offsetQ_1 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1948) begin
                  offsetQ_1 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1948) begin
                    offsetQ_1 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1948) begin
                      offsetQ_1 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1948) begin
                        offsetQ_1 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1948) begin
                          offsetQ_1 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1948) begin
                            offsetQ_1 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1948) begin
                              offsetQ_1 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1948) begin
                                offsetQ_1 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1948) begin
                                  offsetQ_1 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1948) begin
                                    offsetQ_1 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1948) begin
                                      offsetQ_1 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_1 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_2 <= 4'h0;
    end else begin
      if (initBits_2) begin
        if (4'hf == _T_1966) begin
          offsetQ_2 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1966) begin
            offsetQ_2 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1966) begin
              offsetQ_2 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1966) begin
                offsetQ_2 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1966) begin
                  offsetQ_2 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1966) begin
                    offsetQ_2 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1966) begin
                      offsetQ_2 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1966) begin
                        offsetQ_2 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1966) begin
                          offsetQ_2 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1966) begin
                            offsetQ_2 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1966) begin
                              offsetQ_2 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1966) begin
                                offsetQ_2 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1966) begin
                                  offsetQ_2 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1966) begin
                                    offsetQ_2 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1966) begin
                                      offsetQ_2 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_2 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_3 <= 4'h0;
    end else begin
      if (initBits_3) begin
        if (4'hf == _T_1984) begin
          offsetQ_3 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_1984) begin
            offsetQ_3 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_1984) begin
              offsetQ_3 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_1984) begin
                offsetQ_3 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_1984) begin
                  offsetQ_3 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_1984) begin
                    offsetQ_3 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_1984) begin
                      offsetQ_3 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_1984) begin
                        offsetQ_3 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_1984) begin
                          offsetQ_3 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_1984) begin
                            offsetQ_3 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_1984) begin
                              offsetQ_3 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_1984) begin
                                offsetQ_3 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_1984) begin
                                  offsetQ_3 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_1984) begin
                                    offsetQ_3 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_1984) begin
                                      offsetQ_3 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_3 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_4 <= 4'h0;
    end else begin
      if (initBits_4) begin
        if (4'hf == _T_2002) begin
          offsetQ_4 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2002) begin
            offsetQ_4 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2002) begin
              offsetQ_4 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2002) begin
                offsetQ_4 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2002) begin
                  offsetQ_4 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2002) begin
                    offsetQ_4 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2002) begin
                      offsetQ_4 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2002) begin
                        offsetQ_4 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2002) begin
                          offsetQ_4 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2002) begin
                            offsetQ_4 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2002) begin
                              offsetQ_4 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2002) begin
                                offsetQ_4 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2002) begin
                                  offsetQ_4 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2002) begin
                                    offsetQ_4 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2002) begin
                                      offsetQ_4 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_4 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_5 <= 4'h0;
    end else begin
      if (initBits_5) begin
        if (4'hf == _T_2020) begin
          offsetQ_5 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2020) begin
            offsetQ_5 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2020) begin
              offsetQ_5 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2020) begin
                offsetQ_5 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2020) begin
                  offsetQ_5 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2020) begin
                    offsetQ_5 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2020) begin
                      offsetQ_5 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2020) begin
                        offsetQ_5 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2020) begin
                          offsetQ_5 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2020) begin
                            offsetQ_5 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2020) begin
                              offsetQ_5 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2020) begin
                                offsetQ_5 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2020) begin
                                  offsetQ_5 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2020) begin
                                    offsetQ_5 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2020) begin
                                      offsetQ_5 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_5 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_6 <= 4'h0;
    end else begin
      if (initBits_6) begin
        if (4'hf == _T_2038) begin
          offsetQ_6 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2038) begin
            offsetQ_6 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2038) begin
              offsetQ_6 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2038) begin
                offsetQ_6 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2038) begin
                  offsetQ_6 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2038) begin
                    offsetQ_6 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2038) begin
                      offsetQ_6 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2038) begin
                        offsetQ_6 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2038) begin
                          offsetQ_6 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2038) begin
                            offsetQ_6 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2038) begin
                              offsetQ_6 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2038) begin
                                offsetQ_6 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2038) begin
                                  offsetQ_6 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2038) begin
                                    offsetQ_6 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2038) begin
                                      offsetQ_6 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_6 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_7 <= 4'h0;
    end else begin
      if (initBits_7) begin
        if (4'hf == _T_2056) begin
          offsetQ_7 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2056) begin
            offsetQ_7 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2056) begin
              offsetQ_7 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2056) begin
                offsetQ_7 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2056) begin
                  offsetQ_7 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2056) begin
                    offsetQ_7 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2056) begin
                      offsetQ_7 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2056) begin
                        offsetQ_7 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2056) begin
                          offsetQ_7 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2056) begin
                            offsetQ_7 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2056) begin
                              offsetQ_7 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2056) begin
                                offsetQ_7 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2056) begin
                                  offsetQ_7 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2056) begin
                                    offsetQ_7 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2056) begin
                                      offsetQ_7 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_7 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_8 <= 4'h0;
    end else begin
      if (initBits_8) begin
        if (4'hf == _T_2074) begin
          offsetQ_8 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2074) begin
            offsetQ_8 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2074) begin
              offsetQ_8 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2074) begin
                offsetQ_8 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2074) begin
                  offsetQ_8 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2074) begin
                    offsetQ_8 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2074) begin
                      offsetQ_8 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2074) begin
                        offsetQ_8 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2074) begin
                          offsetQ_8 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2074) begin
                            offsetQ_8 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2074) begin
                              offsetQ_8 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2074) begin
                                offsetQ_8 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2074) begin
                                  offsetQ_8 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2074) begin
                                    offsetQ_8 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2074) begin
                                      offsetQ_8 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_8 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_9 <= 4'h0;
    end else begin
      if (initBits_9) begin
        if (4'hf == _T_2092) begin
          offsetQ_9 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2092) begin
            offsetQ_9 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2092) begin
              offsetQ_9 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2092) begin
                offsetQ_9 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2092) begin
                  offsetQ_9 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2092) begin
                    offsetQ_9 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2092) begin
                      offsetQ_9 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2092) begin
                        offsetQ_9 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2092) begin
                          offsetQ_9 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2092) begin
                            offsetQ_9 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2092) begin
                              offsetQ_9 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2092) begin
                                offsetQ_9 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2092) begin
                                  offsetQ_9 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2092) begin
                                    offsetQ_9 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2092) begin
                                      offsetQ_9 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_9 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_10 <= 4'h0;
    end else begin
      if (initBits_10) begin
        if (4'hf == _T_2110) begin
          offsetQ_10 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2110) begin
            offsetQ_10 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2110) begin
              offsetQ_10 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2110) begin
                offsetQ_10 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2110) begin
                  offsetQ_10 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2110) begin
                    offsetQ_10 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2110) begin
                      offsetQ_10 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2110) begin
                        offsetQ_10 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2110) begin
                          offsetQ_10 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2110) begin
                            offsetQ_10 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2110) begin
                              offsetQ_10 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2110) begin
                                offsetQ_10 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2110) begin
                                  offsetQ_10 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2110) begin
                                    offsetQ_10 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2110) begin
                                      offsetQ_10 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_10 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_11 <= 4'h0;
    end else begin
      if (initBits_11) begin
        if (4'hf == _T_2128) begin
          offsetQ_11 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2128) begin
            offsetQ_11 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2128) begin
              offsetQ_11 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2128) begin
                offsetQ_11 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2128) begin
                  offsetQ_11 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2128) begin
                    offsetQ_11 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2128) begin
                      offsetQ_11 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2128) begin
                        offsetQ_11 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2128) begin
                          offsetQ_11 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2128) begin
                            offsetQ_11 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2128) begin
                              offsetQ_11 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2128) begin
                                offsetQ_11 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2128) begin
                                  offsetQ_11 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2128) begin
                                    offsetQ_11 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2128) begin
                                      offsetQ_11 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_11 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_12 <= 4'h0;
    end else begin
      if (initBits_12) begin
        if (4'hf == _T_2146) begin
          offsetQ_12 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2146) begin
            offsetQ_12 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2146) begin
              offsetQ_12 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2146) begin
                offsetQ_12 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2146) begin
                  offsetQ_12 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2146) begin
                    offsetQ_12 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2146) begin
                      offsetQ_12 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2146) begin
                        offsetQ_12 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2146) begin
                          offsetQ_12 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2146) begin
                            offsetQ_12 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2146) begin
                              offsetQ_12 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2146) begin
                                offsetQ_12 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2146) begin
                                  offsetQ_12 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2146) begin
                                    offsetQ_12 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2146) begin
                                      offsetQ_12 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_12 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_13 <= 4'h0;
    end else begin
      if (initBits_13) begin
        if (4'hf == _T_2164) begin
          offsetQ_13 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2164) begin
            offsetQ_13 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2164) begin
              offsetQ_13 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2164) begin
                offsetQ_13 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2164) begin
                  offsetQ_13 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2164) begin
                    offsetQ_13 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2164) begin
                      offsetQ_13 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2164) begin
                        offsetQ_13 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2164) begin
                          offsetQ_13 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2164) begin
                            offsetQ_13 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2164) begin
                              offsetQ_13 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2164) begin
                                offsetQ_13 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2164) begin
                                  offsetQ_13 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2164) begin
                                    offsetQ_13 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2164) begin
                                      offsetQ_13 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_13 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_14 <= 4'h0;
    end else begin
      if (initBits_14) begin
        if (4'hf == _T_2182) begin
          offsetQ_14 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2182) begin
            offsetQ_14 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2182) begin
              offsetQ_14 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2182) begin
                offsetQ_14 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2182) begin
                  offsetQ_14 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2182) begin
                    offsetQ_14 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2182) begin
                      offsetQ_14 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2182) begin
                        offsetQ_14 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2182) begin
                          offsetQ_14 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2182) begin
                            offsetQ_14 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2182) begin
                              offsetQ_14 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2182) begin
                                offsetQ_14 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2182) begin
                                  offsetQ_14 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2182) begin
                                    offsetQ_14 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2182) begin
                                      offsetQ_14 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_14 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      offsetQ_15 <= 4'h0;
    end else begin
      if (initBits_15) begin
        if (4'hf == _T_2200) begin
          offsetQ_15 <= io_bbLoadOffsets_15;
        end else begin
          if (4'he == _T_2200) begin
            offsetQ_15 <= io_bbLoadOffsets_14;
          end else begin
            if (4'hd == _T_2200) begin
              offsetQ_15 <= io_bbLoadOffsets_13;
            end else begin
              if (4'hc == _T_2200) begin
                offsetQ_15 <= io_bbLoadOffsets_12;
              end else begin
                if (4'hb == _T_2200) begin
                  offsetQ_15 <= io_bbLoadOffsets_11;
                end else begin
                  if (4'ha == _T_2200) begin
                    offsetQ_15 <= io_bbLoadOffsets_10;
                  end else begin
                    if (4'h9 == _T_2200) begin
                      offsetQ_15 <= io_bbLoadOffsets_9;
                    end else begin
                      if (4'h8 == _T_2200) begin
                        offsetQ_15 <= io_bbLoadOffsets_8;
                      end else begin
                        if (4'h7 == _T_2200) begin
                          offsetQ_15 <= io_bbLoadOffsets_7;
                        end else begin
                          if (4'h6 == _T_2200) begin
                            offsetQ_15 <= io_bbLoadOffsets_6;
                          end else begin
                            if (4'h5 == _T_2200) begin
                              offsetQ_15 <= io_bbLoadOffsets_5;
                            end else begin
                              if (4'h4 == _T_2200) begin
                                offsetQ_15 <= io_bbLoadOffsets_4;
                              end else begin
                                if (4'h3 == _T_2200) begin
                                  offsetQ_15 <= io_bbLoadOffsets_3;
                                end else begin
                                  if (4'h2 == _T_2200) begin
                                    offsetQ_15 <= io_bbLoadOffsets_2;
                                  end else begin
                                    if (4'h1 == _T_2200) begin
                                      offsetQ_15 <= io_bbLoadOffsets_1;
                                    end else begin
                                      offsetQ_15 <= io_bbLoadOffsets_0;
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      portQ_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        portQ_0 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        portQ_1 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        portQ_2 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        portQ_3 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        portQ_4 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        portQ_5 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        portQ_6 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        portQ_7 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        portQ_8 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        portQ_9 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        portQ_10 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        portQ_11 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        portQ_12 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        portQ_13 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        portQ_14 <= 1'h0;
      end
    end
    if (reset) begin
      portQ_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        portQ_15 <= 1'h0;
      end
    end
    if (reset) begin
      addrQ_0 <= 31'h0;
    end else begin
      if (!(initBits_0)) begin
        if (_T_97704) begin
          addrQ_0 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_1 <= 31'h0;
    end else begin
      if (!(initBits_1)) begin
        if (_T_97719) begin
          addrQ_1 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_2 <= 31'h0;
    end else begin
      if (!(initBits_2)) begin
        if (_T_97734) begin
          addrQ_2 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_3 <= 31'h0;
    end else begin
      if (!(initBits_3)) begin
        if (_T_97749) begin
          addrQ_3 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_4 <= 31'h0;
    end else begin
      if (!(initBits_4)) begin
        if (_T_97764) begin
          addrQ_4 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_5 <= 31'h0;
    end else begin
      if (!(initBits_5)) begin
        if (_T_97779) begin
          addrQ_5 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_6 <= 31'h0;
    end else begin
      if (!(initBits_6)) begin
        if (_T_97794) begin
          addrQ_6 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_7 <= 31'h0;
    end else begin
      if (!(initBits_7)) begin
        if (_T_97809) begin
          addrQ_7 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_8 <= 31'h0;
    end else begin
      if (!(initBits_8)) begin
        if (_T_97824) begin
          addrQ_8 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_9 <= 31'h0;
    end else begin
      if (!(initBits_9)) begin
        if (_T_97839) begin
          addrQ_9 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_10 <= 31'h0;
    end else begin
      if (!(initBits_10)) begin
        if (_T_97854) begin
          addrQ_10 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_11 <= 31'h0;
    end else begin
      if (!(initBits_11)) begin
        if (_T_97869) begin
          addrQ_11 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_12 <= 31'h0;
    end else begin
      if (!(initBits_12)) begin
        if (_T_97884) begin
          addrQ_12 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_13 <= 31'h0;
    end else begin
      if (!(initBits_13)) begin
        if (_T_97899) begin
          addrQ_13 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_14 <= 31'h0;
    end else begin
      if (!(initBits_14)) begin
        if (_T_97914) begin
          addrQ_14 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      addrQ_15 <= 31'h0;
    end else begin
      if (!(initBits_15)) begin
        if (_T_97929) begin
          addrQ_15 <= io_addrFromLoadPorts_0;
        end
      end
    end
    if (reset) begin
      dataQ_0 <= 32'h0;
    end else begin
      if (bypassRequest_0) begin
        if (_T_88304) begin
          if (4'hf == _T_88287) begin
            dataQ_0 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88287) begin
              dataQ_0 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88287) begin
                dataQ_0 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88287) begin
                  dataQ_0 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88287) begin
                    dataQ_0 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88287) begin
                      dataQ_0 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88287) begin
                        dataQ_0 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88287) begin
                          dataQ_0 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88287) begin
                            dataQ_0 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88287) begin
                              dataQ_0 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88287) begin
                                dataQ_0 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88287) begin
                                  dataQ_0 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88287) begin
                                    dataQ_0 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88287) begin
                                      dataQ_0 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88287) begin
                                        dataQ_0 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_0 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_0 <= 32'h0;
        end
      end else begin
        if (_T_93694) begin
          dataQ_0 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_1 <= 32'h0;
    end else begin
      if (bypassRequest_1) begin
        if (_T_88440) begin
          if (4'hf == _T_88423) begin
            dataQ_1 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88423) begin
              dataQ_1 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88423) begin
                dataQ_1 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88423) begin
                  dataQ_1 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88423) begin
                    dataQ_1 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88423) begin
                      dataQ_1 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88423) begin
                        dataQ_1 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88423) begin
                          dataQ_1 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88423) begin
                            dataQ_1 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88423) begin
                              dataQ_1 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88423) begin
                                dataQ_1 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88423) begin
                                  dataQ_1 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88423) begin
                                    dataQ_1 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88423) begin
                                      dataQ_1 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88423) begin
                                        dataQ_1 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_1 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_1 <= 32'h0;
        end
      end else begin
        if (_T_93700) begin
          dataQ_1 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_2 <= 32'h0;
    end else begin
      if (bypassRequest_2) begin
        if (_T_88576) begin
          if (4'hf == _T_88559) begin
            dataQ_2 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88559) begin
              dataQ_2 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88559) begin
                dataQ_2 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88559) begin
                  dataQ_2 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88559) begin
                    dataQ_2 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88559) begin
                      dataQ_2 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88559) begin
                        dataQ_2 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88559) begin
                          dataQ_2 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88559) begin
                            dataQ_2 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88559) begin
                              dataQ_2 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88559) begin
                                dataQ_2 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88559) begin
                                  dataQ_2 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88559) begin
                                    dataQ_2 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88559) begin
                                      dataQ_2 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88559) begin
                                        dataQ_2 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_2 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_2 <= 32'h0;
        end
      end else begin
        if (_T_93706) begin
          dataQ_2 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_3 <= 32'h0;
    end else begin
      if (bypassRequest_3) begin
        if (_T_88712) begin
          if (4'hf == _T_88695) begin
            dataQ_3 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88695) begin
              dataQ_3 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88695) begin
                dataQ_3 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88695) begin
                  dataQ_3 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88695) begin
                    dataQ_3 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88695) begin
                      dataQ_3 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88695) begin
                        dataQ_3 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88695) begin
                          dataQ_3 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88695) begin
                            dataQ_3 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88695) begin
                              dataQ_3 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88695) begin
                                dataQ_3 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88695) begin
                                  dataQ_3 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88695) begin
                                    dataQ_3 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88695) begin
                                      dataQ_3 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88695) begin
                                        dataQ_3 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_3 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_3 <= 32'h0;
        end
      end else begin
        if (_T_93712) begin
          dataQ_3 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_4 <= 32'h0;
    end else begin
      if (bypassRequest_4) begin
        if (_T_88848) begin
          if (4'hf == _T_88831) begin
            dataQ_4 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88831) begin
              dataQ_4 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88831) begin
                dataQ_4 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88831) begin
                  dataQ_4 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88831) begin
                    dataQ_4 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88831) begin
                      dataQ_4 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88831) begin
                        dataQ_4 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88831) begin
                          dataQ_4 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88831) begin
                            dataQ_4 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88831) begin
                              dataQ_4 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88831) begin
                                dataQ_4 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88831) begin
                                  dataQ_4 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88831) begin
                                    dataQ_4 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88831) begin
                                      dataQ_4 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88831) begin
                                        dataQ_4 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_4 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_4 <= 32'h0;
        end
      end else begin
        if (_T_93718) begin
          dataQ_4 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_5 <= 32'h0;
    end else begin
      if (bypassRequest_5) begin
        if (_T_88984) begin
          if (4'hf == _T_88967) begin
            dataQ_5 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_88967) begin
              dataQ_5 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_88967) begin
                dataQ_5 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_88967) begin
                  dataQ_5 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_88967) begin
                    dataQ_5 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_88967) begin
                      dataQ_5 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_88967) begin
                        dataQ_5 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_88967) begin
                          dataQ_5 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_88967) begin
                            dataQ_5 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_88967) begin
                              dataQ_5 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_88967) begin
                                dataQ_5 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_88967) begin
                                  dataQ_5 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_88967) begin
                                    dataQ_5 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_88967) begin
                                      dataQ_5 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_88967) begin
                                        dataQ_5 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_5 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_5 <= 32'h0;
        end
      end else begin
        if (_T_93724) begin
          dataQ_5 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_6 <= 32'h0;
    end else begin
      if (bypassRequest_6) begin
        if (_T_89120) begin
          if (4'hf == _T_89103) begin
            dataQ_6 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89103) begin
              dataQ_6 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89103) begin
                dataQ_6 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89103) begin
                  dataQ_6 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89103) begin
                    dataQ_6 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89103) begin
                      dataQ_6 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89103) begin
                        dataQ_6 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89103) begin
                          dataQ_6 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89103) begin
                            dataQ_6 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89103) begin
                              dataQ_6 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89103) begin
                                dataQ_6 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89103) begin
                                  dataQ_6 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89103) begin
                                    dataQ_6 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89103) begin
                                      dataQ_6 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89103) begin
                                        dataQ_6 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_6 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_6 <= 32'h0;
        end
      end else begin
        if (_T_93730) begin
          dataQ_6 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_7 <= 32'h0;
    end else begin
      if (bypassRequest_7) begin
        if (_T_89256) begin
          if (4'hf == _T_89239) begin
            dataQ_7 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89239) begin
              dataQ_7 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89239) begin
                dataQ_7 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89239) begin
                  dataQ_7 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89239) begin
                    dataQ_7 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89239) begin
                      dataQ_7 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89239) begin
                        dataQ_7 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89239) begin
                          dataQ_7 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89239) begin
                            dataQ_7 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89239) begin
                              dataQ_7 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89239) begin
                                dataQ_7 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89239) begin
                                  dataQ_7 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89239) begin
                                    dataQ_7 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89239) begin
                                      dataQ_7 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89239) begin
                                        dataQ_7 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_7 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_7 <= 32'h0;
        end
      end else begin
        if (_T_93736) begin
          dataQ_7 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_8 <= 32'h0;
    end else begin
      if (bypassRequest_8) begin
        if (_T_89392) begin
          if (4'hf == _T_89375) begin
            dataQ_8 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89375) begin
              dataQ_8 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89375) begin
                dataQ_8 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89375) begin
                  dataQ_8 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89375) begin
                    dataQ_8 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89375) begin
                      dataQ_8 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89375) begin
                        dataQ_8 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89375) begin
                          dataQ_8 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89375) begin
                            dataQ_8 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89375) begin
                              dataQ_8 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89375) begin
                                dataQ_8 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89375) begin
                                  dataQ_8 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89375) begin
                                    dataQ_8 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89375) begin
                                      dataQ_8 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89375) begin
                                        dataQ_8 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_8 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_8 <= 32'h0;
        end
      end else begin
        if (_T_93742) begin
          dataQ_8 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_9 <= 32'h0;
    end else begin
      if (bypassRequest_9) begin
        if (_T_89528) begin
          if (4'hf == _T_89511) begin
            dataQ_9 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89511) begin
              dataQ_9 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89511) begin
                dataQ_9 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89511) begin
                  dataQ_9 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89511) begin
                    dataQ_9 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89511) begin
                      dataQ_9 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89511) begin
                        dataQ_9 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89511) begin
                          dataQ_9 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89511) begin
                            dataQ_9 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89511) begin
                              dataQ_9 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89511) begin
                                dataQ_9 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89511) begin
                                  dataQ_9 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89511) begin
                                    dataQ_9 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89511) begin
                                      dataQ_9 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89511) begin
                                        dataQ_9 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_9 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_9 <= 32'h0;
        end
      end else begin
        if (_T_93748) begin
          dataQ_9 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_10 <= 32'h0;
    end else begin
      if (bypassRequest_10) begin
        if (_T_89664) begin
          if (4'hf == _T_89647) begin
            dataQ_10 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89647) begin
              dataQ_10 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89647) begin
                dataQ_10 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89647) begin
                  dataQ_10 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89647) begin
                    dataQ_10 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89647) begin
                      dataQ_10 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89647) begin
                        dataQ_10 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89647) begin
                          dataQ_10 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89647) begin
                            dataQ_10 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89647) begin
                              dataQ_10 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89647) begin
                                dataQ_10 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89647) begin
                                  dataQ_10 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89647) begin
                                    dataQ_10 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89647) begin
                                      dataQ_10 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89647) begin
                                        dataQ_10 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_10 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_10 <= 32'h0;
        end
      end else begin
        if (_T_93754) begin
          dataQ_10 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_11 <= 32'h0;
    end else begin
      if (bypassRequest_11) begin
        if (_T_89800) begin
          if (4'hf == _T_89783) begin
            dataQ_11 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89783) begin
              dataQ_11 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89783) begin
                dataQ_11 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89783) begin
                  dataQ_11 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89783) begin
                    dataQ_11 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89783) begin
                      dataQ_11 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89783) begin
                        dataQ_11 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89783) begin
                          dataQ_11 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89783) begin
                            dataQ_11 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89783) begin
                              dataQ_11 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89783) begin
                                dataQ_11 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89783) begin
                                  dataQ_11 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89783) begin
                                    dataQ_11 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89783) begin
                                      dataQ_11 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89783) begin
                                        dataQ_11 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_11 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_11 <= 32'h0;
        end
      end else begin
        if (_T_93760) begin
          dataQ_11 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_12 <= 32'h0;
    end else begin
      if (bypassRequest_12) begin
        if (_T_89936) begin
          if (4'hf == _T_89919) begin
            dataQ_12 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_89919) begin
              dataQ_12 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_89919) begin
                dataQ_12 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_89919) begin
                  dataQ_12 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_89919) begin
                    dataQ_12 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_89919) begin
                      dataQ_12 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_89919) begin
                        dataQ_12 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_89919) begin
                          dataQ_12 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_89919) begin
                            dataQ_12 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_89919) begin
                              dataQ_12 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_89919) begin
                                dataQ_12 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_89919) begin
                                  dataQ_12 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_89919) begin
                                    dataQ_12 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_89919) begin
                                      dataQ_12 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_89919) begin
                                        dataQ_12 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_12 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_12 <= 32'h0;
        end
      end else begin
        if (_T_93766) begin
          dataQ_12 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_13 <= 32'h0;
    end else begin
      if (bypassRequest_13) begin
        if (_T_90072) begin
          if (4'hf == _T_90055) begin
            dataQ_13 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90055) begin
              dataQ_13 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90055) begin
                dataQ_13 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90055) begin
                  dataQ_13 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90055) begin
                    dataQ_13 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90055) begin
                      dataQ_13 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90055) begin
                        dataQ_13 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90055) begin
                          dataQ_13 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90055) begin
                            dataQ_13 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90055) begin
                              dataQ_13 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90055) begin
                                dataQ_13 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90055) begin
                                  dataQ_13 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90055) begin
                                    dataQ_13 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90055) begin
                                      dataQ_13 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90055) begin
                                        dataQ_13 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_13 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_13 <= 32'h0;
        end
      end else begin
        if (_T_93772) begin
          dataQ_13 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_14 <= 32'h0;
    end else begin
      if (bypassRequest_14) begin
        if (_T_90208) begin
          if (4'hf == _T_90191) begin
            dataQ_14 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90191) begin
              dataQ_14 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90191) begin
                dataQ_14 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90191) begin
                  dataQ_14 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90191) begin
                    dataQ_14 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90191) begin
                      dataQ_14 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90191) begin
                        dataQ_14 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90191) begin
                          dataQ_14 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90191) begin
                            dataQ_14 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90191) begin
                              dataQ_14 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90191) begin
                                dataQ_14 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90191) begin
                                  dataQ_14 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90191) begin
                                    dataQ_14 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90191) begin
                                      dataQ_14 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90191) begin
                                        dataQ_14 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_14 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_14 <= 32'h0;
        end
      end else begin
        if (_T_93778) begin
          dataQ_14 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      dataQ_15 <= 32'h0;
    end else begin
      if (bypassRequest_15) begin
        if (_T_90344) begin
          if (4'hf == _T_90327) begin
            dataQ_15 <= shiftedStoreDataQPreg_15;
          end else begin
            if (4'he == _T_90327) begin
              dataQ_15 <= shiftedStoreDataQPreg_14;
            end else begin
              if (4'hd == _T_90327) begin
                dataQ_15 <= shiftedStoreDataQPreg_13;
              end else begin
                if (4'hc == _T_90327) begin
                  dataQ_15 <= shiftedStoreDataQPreg_12;
                end else begin
                  if (4'hb == _T_90327) begin
                    dataQ_15 <= shiftedStoreDataQPreg_11;
                  end else begin
                    if (4'ha == _T_90327) begin
                      dataQ_15 <= shiftedStoreDataQPreg_10;
                    end else begin
                      if (4'h9 == _T_90327) begin
                        dataQ_15 <= shiftedStoreDataQPreg_9;
                      end else begin
                        if (4'h8 == _T_90327) begin
                          dataQ_15 <= shiftedStoreDataQPreg_8;
                        end else begin
                          if (4'h7 == _T_90327) begin
                            dataQ_15 <= shiftedStoreDataQPreg_7;
                          end else begin
                            if (4'h6 == _T_90327) begin
                              dataQ_15 <= shiftedStoreDataQPreg_6;
                            end else begin
                              if (4'h5 == _T_90327) begin
                                dataQ_15 <= shiftedStoreDataQPreg_5;
                              end else begin
                                if (4'h4 == _T_90327) begin
                                  dataQ_15 <= shiftedStoreDataQPreg_4;
                                end else begin
                                  if (4'h3 == _T_90327) begin
                                    dataQ_15 <= shiftedStoreDataQPreg_3;
                                  end else begin
                                    if (4'h2 == _T_90327) begin
                                      dataQ_15 <= shiftedStoreDataQPreg_2;
                                    end else begin
                                      if (4'h1 == _T_90327) begin
                                        dataQ_15 <= shiftedStoreDataQPreg_1;
                                      end else begin
                                        dataQ_15 <= shiftedStoreDataQPreg_0;
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          dataQ_15 <= 32'h0;
        end
      end else begin
        if (_T_93784) begin
          dataQ_15 <= io_loadDataFromMem;
        end
      end
    end
    if (reset) begin
      addrKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        addrKnown_0 <= 1'h0;
      end else begin
        if (_T_97704) begin
          addrKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        addrKnown_1 <= 1'h0;
      end else begin
        if (_T_97719) begin
          addrKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        addrKnown_2 <= 1'h0;
      end else begin
        if (_T_97734) begin
          addrKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        addrKnown_3 <= 1'h0;
      end else begin
        if (_T_97749) begin
          addrKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        addrKnown_4 <= 1'h0;
      end else begin
        if (_T_97764) begin
          addrKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        addrKnown_5 <= 1'h0;
      end else begin
        if (_T_97779) begin
          addrKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        addrKnown_6 <= 1'h0;
      end else begin
        if (_T_97794) begin
          addrKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        addrKnown_7 <= 1'h0;
      end else begin
        if (_T_97809) begin
          addrKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        addrKnown_8 <= 1'h0;
      end else begin
        if (_T_97824) begin
          addrKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        addrKnown_9 <= 1'h0;
      end else begin
        if (_T_97839) begin
          addrKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        addrKnown_10 <= 1'h0;
      end else begin
        if (_T_97854) begin
          addrKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        addrKnown_11 <= 1'h0;
      end else begin
        if (_T_97869) begin
          addrKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        addrKnown_12 <= 1'h0;
      end else begin
        if (_T_97884) begin
          addrKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        addrKnown_13 <= 1'h0;
      end else begin
        if (_T_97899) begin
          addrKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        addrKnown_14 <= 1'h0;
      end else begin
        if (_T_97914) begin
          addrKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      addrKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        addrKnown_15 <= 1'h0;
      end else begin
        if (_T_97929) begin
          addrKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        dataKnown_0 <= 1'h0;
      end else begin
        if (_T_93695) begin
          dataKnown_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        dataKnown_1 <= 1'h0;
      end else begin
        if (_T_93701) begin
          dataKnown_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        dataKnown_2 <= 1'h0;
      end else begin
        if (_T_93707) begin
          dataKnown_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        dataKnown_3 <= 1'h0;
      end else begin
        if (_T_93713) begin
          dataKnown_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        dataKnown_4 <= 1'h0;
      end else begin
        if (_T_93719) begin
          dataKnown_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        dataKnown_5 <= 1'h0;
      end else begin
        if (_T_93725) begin
          dataKnown_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        dataKnown_6 <= 1'h0;
      end else begin
        if (_T_93731) begin
          dataKnown_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        dataKnown_7 <= 1'h0;
      end else begin
        if (_T_93737) begin
          dataKnown_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        dataKnown_8 <= 1'h0;
      end else begin
        if (_T_93743) begin
          dataKnown_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        dataKnown_9 <= 1'h0;
      end else begin
        if (_T_93749) begin
          dataKnown_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        dataKnown_10 <= 1'h0;
      end else begin
        if (_T_93755) begin
          dataKnown_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        dataKnown_11 <= 1'h0;
      end else begin
        if (_T_93761) begin
          dataKnown_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        dataKnown_12 <= 1'h0;
      end else begin
        if (_T_93767) begin
          dataKnown_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        dataKnown_13 <= 1'h0;
      end else begin
        if (_T_93773) begin
          dataKnown_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        dataKnown_14 <= 1'h0;
      end else begin
        if (_T_93779) begin
          dataKnown_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      dataKnown_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        dataKnown_15 <= 1'h0;
      end else begin
        if (_T_93785) begin
          dataKnown_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        loadCompleted_0 <= 1'h0;
      end else begin
        if (loadCompleting_0) begin
          loadCompleted_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        loadCompleted_1 <= 1'h0;
      end else begin
        if (loadCompleting_1) begin
          loadCompleted_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        loadCompleted_2 <= 1'h0;
      end else begin
        if (loadCompleting_2) begin
          loadCompleted_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        loadCompleted_3 <= 1'h0;
      end else begin
        if (loadCompleting_3) begin
          loadCompleted_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        loadCompleted_4 <= 1'h0;
      end else begin
        if (loadCompleting_4) begin
          loadCompleted_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        loadCompleted_5 <= 1'h0;
      end else begin
        if (loadCompleting_5) begin
          loadCompleted_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        loadCompleted_6 <= 1'h0;
      end else begin
        if (loadCompleting_6) begin
          loadCompleted_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        loadCompleted_7 <= 1'h0;
      end else begin
        if (loadCompleting_7) begin
          loadCompleted_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        loadCompleted_8 <= 1'h0;
      end else begin
        if (loadCompleting_8) begin
          loadCompleted_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        loadCompleted_9 <= 1'h0;
      end else begin
        if (loadCompleting_9) begin
          loadCompleted_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        loadCompleted_10 <= 1'h0;
      end else begin
        if (loadCompleting_10) begin
          loadCompleted_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        loadCompleted_11 <= 1'h0;
      end else begin
        if (loadCompleting_11) begin
          loadCompleted_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        loadCompleted_12 <= 1'h0;
      end else begin
        if (loadCompleting_12) begin
          loadCompleted_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        loadCompleted_13 <= 1'h0;
      end else begin
        if (loadCompleting_13) begin
          loadCompleted_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        loadCompleted_14 <= 1'h0;
      end else begin
        if (loadCompleting_14) begin
          loadCompleted_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadCompleted_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        loadCompleted_15 <= 1'h0;
      end else begin
        if (loadCompleting_15) begin
          loadCompleted_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      allocatedEntries_0 <= 1'h0;
    end else begin
      allocatedEntries_0 <= _T_1884;
    end
    if (reset) begin
      allocatedEntries_1 <= 1'h0;
    end else begin
      allocatedEntries_1 <= _T_1885;
    end
    if (reset) begin
      allocatedEntries_2 <= 1'h0;
    end else begin
      allocatedEntries_2 <= _T_1886;
    end
    if (reset) begin
      allocatedEntries_3 <= 1'h0;
    end else begin
      allocatedEntries_3 <= _T_1887;
    end
    if (reset) begin
      allocatedEntries_4 <= 1'h0;
    end else begin
      allocatedEntries_4 <= _T_1888;
    end
    if (reset) begin
      allocatedEntries_5 <= 1'h0;
    end else begin
      allocatedEntries_5 <= _T_1889;
    end
    if (reset) begin
      allocatedEntries_6 <= 1'h0;
    end else begin
      allocatedEntries_6 <= _T_1890;
    end
    if (reset) begin
      allocatedEntries_7 <= 1'h0;
    end else begin
      allocatedEntries_7 <= _T_1891;
    end
    if (reset) begin
      allocatedEntries_8 <= 1'h0;
    end else begin
      allocatedEntries_8 <= _T_1892;
    end
    if (reset) begin
      allocatedEntries_9 <= 1'h0;
    end else begin
      allocatedEntries_9 <= _T_1893;
    end
    if (reset) begin
      allocatedEntries_10 <= 1'h0;
    end else begin
      allocatedEntries_10 <= _T_1894;
    end
    if (reset) begin
      allocatedEntries_11 <= 1'h0;
    end else begin
      allocatedEntries_11 <= _T_1895;
    end
    if (reset) begin
      allocatedEntries_12 <= 1'h0;
    end else begin
      allocatedEntries_12 <= _T_1896;
    end
    if (reset) begin
      allocatedEntries_13 <= 1'h0;
    end else begin
      allocatedEntries_13 <= _T_1897;
    end
    if (reset) begin
      allocatedEntries_14 <= 1'h0;
    end else begin
      allocatedEntries_14 <= _T_1898;
    end
    if (reset) begin
      allocatedEntries_15 <= 1'h0;
    end else begin
      allocatedEntries_15 <= _T_1899;
    end
    if (reset) begin
      bypassInitiated_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        bypassInitiated_0 <= 1'h0;
      end else begin
        if (bypassRequest_0) begin
          bypassInitiated_0 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        bypassInitiated_1 <= 1'h0;
      end else begin
        if (bypassRequest_1) begin
          bypassInitiated_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        bypassInitiated_2 <= 1'h0;
      end else begin
        if (bypassRequest_2) begin
          bypassInitiated_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        bypassInitiated_3 <= 1'h0;
      end else begin
        if (bypassRequest_3) begin
          bypassInitiated_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        bypassInitiated_4 <= 1'h0;
      end else begin
        if (bypassRequest_4) begin
          bypassInitiated_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        bypassInitiated_5 <= 1'h0;
      end else begin
        if (bypassRequest_5) begin
          bypassInitiated_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        bypassInitiated_6 <= 1'h0;
      end else begin
        if (bypassRequest_6) begin
          bypassInitiated_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        bypassInitiated_7 <= 1'h0;
      end else begin
        if (bypassRequest_7) begin
          bypassInitiated_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        bypassInitiated_8 <= 1'h0;
      end else begin
        if (bypassRequest_8) begin
          bypassInitiated_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        bypassInitiated_9 <= 1'h0;
      end else begin
        if (bypassRequest_9) begin
          bypassInitiated_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        bypassInitiated_10 <= 1'h0;
      end else begin
        if (bypassRequest_10) begin
          bypassInitiated_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        bypassInitiated_11 <= 1'h0;
      end else begin
        if (bypassRequest_11) begin
          bypassInitiated_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        bypassInitiated_12 <= 1'h0;
      end else begin
        if (bypassRequest_12) begin
          bypassInitiated_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        bypassInitiated_13 <= 1'h0;
      end else begin
        if (bypassRequest_13) begin
          bypassInitiated_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        bypassInitiated_14 <= 1'h0;
      end else begin
        if (bypassRequest_14) begin
          bypassInitiated_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      bypassInitiated_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        bypassInitiated_15 <= 1'h0;
      end else begin
        if (bypassRequest_15) begin
          bypassInitiated_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      checkBits_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        checkBits_0 <= _T_2227;
      end else begin
        if (io_storeEmpty) begin
          checkBits_0 <= 1'h0;
        end else begin
          if (_T_2231) begin
            checkBits_0 <= 1'h0;
          end else begin
            if (_T_2239) begin
              checkBits_0 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        checkBits_1 <= _T_2257;
      end else begin
        if (io_storeEmpty) begin
          checkBits_1 <= 1'h0;
        end else begin
          if (_T_2261) begin
            checkBits_1 <= 1'h0;
          end else begin
            if (_T_2269) begin
              checkBits_1 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        checkBits_2 <= _T_2287;
      end else begin
        if (io_storeEmpty) begin
          checkBits_2 <= 1'h0;
        end else begin
          if (_T_2291) begin
            checkBits_2 <= 1'h0;
          end else begin
            if (_T_2299) begin
              checkBits_2 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        checkBits_3 <= _T_2317;
      end else begin
        if (io_storeEmpty) begin
          checkBits_3 <= 1'h0;
        end else begin
          if (_T_2321) begin
            checkBits_3 <= 1'h0;
          end else begin
            if (_T_2329) begin
              checkBits_3 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        checkBits_4 <= _T_2347;
      end else begin
        if (io_storeEmpty) begin
          checkBits_4 <= 1'h0;
        end else begin
          if (_T_2351) begin
            checkBits_4 <= 1'h0;
          end else begin
            if (_T_2359) begin
              checkBits_4 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        checkBits_5 <= _T_2377;
      end else begin
        if (io_storeEmpty) begin
          checkBits_5 <= 1'h0;
        end else begin
          if (_T_2381) begin
            checkBits_5 <= 1'h0;
          end else begin
            if (_T_2389) begin
              checkBits_5 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        checkBits_6 <= _T_2407;
      end else begin
        if (io_storeEmpty) begin
          checkBits_6 <= 1'h0;
        end else begin
          if (_T_2411) begin
            checkBits_6 <= 1'h0;
          end else begin
            if (_T_2419) begin
              checkBits_6 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        checkBits_7 <= _T_2437;
      end else begin
        if (io_storeEmpty) begin
          checkBits_7 <= 1'h0;
        end else begin
          if (_T_2441) begin
            checkBits_7 <= 1'h0;
          end else begin
            if (_T_2449) begin
              checkBits_7 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        checkBits_8 <= _T_2467;
      end else begin
        if (io_storeEmpty) begin
          checkBits_8 <= 1'h0;
        end else begin
          if (_T_2471) begin
            checkBits_8 <= 1'h0;
          end else begin
            if (_T_2479) begin
              checkBits_8 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        checkBits_9 <= _T_2497;
      end else begin
        if (io_storeEmpty) begin
          checkBits_9 <= 1'h0;
        end else begin
          if (_T_2501) begin
            checkBits_9 <= 1'h0;
          end else begin
            if (_T_2509) begin
              checkBits_9 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        checkBits_10 <= _T_2527;
      end else begin
        if (io_storeEmpty) begin
          checkBits_10 <= 1'h0;
        end else begin
          if (_T_2531) begin
            checkBits_10 <= 1'h0;
          end else begin
            if (_T_2539) begin
              checkBits_10 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        checkBits_11 <= _T_2557;
      end else begin
        if (io_storeEmpty) begin
          checkBits_11 <= 1'h0;
        end else begin
          if (_T_2561) begin
            checkBits_11 <= 1'h0;
          end else begin
            if (_T_2569) begin
              checkBits_11 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        checkBits_12 <= _T_2587;
      end else begin
        if (io_storeEmpty) begin
          checkBits_12 <= 1'h0;
        end else begin
          if (_T_2591) begin
            checkBits_12 <= 1'h0;
          end else begin
            if (_T_2599) begin
              checkBits_12 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        checkBits_13 <= _T_2617;
      end else begin
        if (io_storeEmpty) begin
          checkBits_13 <= 1'h0;
        end else begin
          if (_T_2621) begin
            checkBits_13 <= 1'h0;
          end else begin
            if (_T_2629) begin
              checkBits_13 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        checkBits_14 <= _T_2647;
      end else begin
        if (io_storeEmpty) begin
          checkBits_14 <= 1'h0;
        end else begin
          if (_T_2651) begin
            checkBits_14 <= 1'h0;
          end else begin
            if (_T_2659) begin
              checkBits_14 <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      checkBits_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        checkBits_15 <= _T_2677;
      end else begin
        if (io_storeEmpty) begin
          checkBits_15 <= 1'h0;
        end else begin
          if (_T_2681) begin
            checkBits_15 <= 1'h0;
          end else begin
            if (_T_2689) begin
              checkBits_15 <= 1'h0;
            end
          end
        end
      end
    end
    previousStoreHead <= io_storeHead;
    conflictPReg_0_0 <= _T_18288[0];
    conflictPReg_0_1 <= _T_18288[1];
    conflictPReg_0_2 <= _T_18288[2];
    conflictPReg_0_3 <= _T_18288[3];
    conflictPReg_0_4 <= _T_18288[4];
    conflictPReg_0_5 <= _T_18288[5];
    conflictPReg_0_6 <= _T_18288[6];
    conflictPReg_0_7 <= _T_18288[7];
    conflictPReg_0_8 <= _T_18288[8];
    conflictPReg_0_9 <= _T_18288[9];
    conflictPReg_0_10 <= _T_18288[10];
    conflictPReg_0_11 <= _T_18288[11];
    conflictPReg_0_12 <= _T_18288[12];
    conflictPReg_0_13 <= _T_18288[13];
    conflictPReg_0_14 <= _T_18288[14];
    conflictPReg_0_15 <= _T_18288[15];
    conflictPReg_1_0 <= _T_19146[0];
    conflictPReg_1_1 <= _T_19146[1];
    conflictPReg_1_2 <= _T_19146[2];
    conflictPReg_1_3 <= _T_19146[3];
    conflictPReg_1_4 <= _T_19146[4];
    conflictPReg_1_5 <= _T_19146[5];
    conflictPReg_1_6 <= _T_19146[6];
    conflictPReg_1_7 <= _T_19146[7];
    conflictPReg_1_8 <= _T_19146[8];
    conflictPReg_1_9 <= _T_19146[9];
    conflictPReg_1_10 <= _T_19146[10];
    conflictPReg_1_11 <= _T_19146[11];
    conflictPReg_1_12 <= _T_19146[12];
    conflictPReg_1_13 <= _T_19146[13];
    conflictPReg_1_14 <= _T_19146[14];
    conflictPReg_1_15 <= _T_19146[15];
    conflictPReg_2_0 <= _T_20004[0];
    conflictPReg_2_1 <= _T_20004[1];
    conflictPReg_2_2 <= _T_20004[2];
    conflictPReg_2_3 <= _T_20004[3];
    conflictPReg_2_4 <= _T_20004[4];
    conflictPReg_2_5 <= _T_20004[5];
    conflictPReg_2_6 <= _T_20004[6];
    conflictPReg_2_7 <= _T_20004[7];
    conflictPReg_2_8 <= _T_20004[8];
    conflictPReg_2_9 <= _T_20004[9];
    conflictPReg_2_10 <= _T_20004[10];
    conflictPReg_2_11 <= _T_20004[11];
    conflictPReg_2_12 <= _T_20004[12];
    conflictPReg_2_13 <= _T_20004[13];
    conflictPReg_2_14 <= _T_20004[14];
    conflictPReg_2_15 <= _T_20004[15];
    conflictPReg_3_0 <= _T_20862[0];
    conflictPReg_3_1 <= _T_20862[1];
    conflictPReg_3_2 <= _T_20862[2];
    conflictPReg_3_3 <= _T_20862[3];
    conflictPReg_3_4 <= _T_20862[4];
    conflictPReg_3_5 <= _T_20862[5];
    conflictPReg_3_6 <= _T_20862[6];
    conflictPReg_3_7 <= _T_20862[7];
    conflictPReg_3_8 <= _T_20862[8];
    conflictPReg_3_9 <= _T_20862[9];
    conflictPReg_3_10 <= _T_20862[10];
    conflictPReg_3_11 <= _T_20862[11];
    conflictPReg_3_12 <= _T_20862[12];
    conflictPReg_3_13 <= _T_20862[13];
    conflictPReg_3_14 <= _T_20862[14];
    conflictPReg_3_15 <= _T_20862[15];
    conflictPReg_4_0 <= _T_21720[0];
    conflictPReg_4_1 <= _T_21720[1];
    conflictPReg_4_2 <= _T_21720[2];
    conflictPReg_4_3 <= _T_21720[3];
    conflictPReg_4_4 <= _T_21720[4];
    conflictPReg_4_5 <= _T_21720[5];
    conflictPReg_4_6 <= _T_21720[6];
    conflictPReg_4_7 <= _T_21720[7];
    conflictPReg_4_8 <= _T_21720[8];
    conflictPReg_4_9 <= _T_21720[9];
    conflictPReg_4_10 <= _T_21720[10];
    conflictPReg_4_11 <= _T_21720[11];
    conflictPReg_4_12 <= _T_21720[12];
    conflictPReg_4_13 <= _T_21720[13];
    conflictPReg_4_14 <= _T_21720[14];
    conflictPReg_4_15 <= _T_21720[15];
    conflictPReg_5_0 <= _T_22578[0];
    conflictPReg_5_1 <= _T_22578[1];
    conflictPReg_5_2 <= _T_22578[2];
    conflictPReg_5_3 <= _T_22578[3];
    conflictPReg_5_4 <= _T_22578[4];
    conflictPReg_5_5 <= _T_22578[5];
    conflictPReg_5_6 <= _T_22578[6];
    conflictPReg_5_7 <= _T_22578[7];
    conflictPReg_5_8 <= _T_22578[8];
    conflictPReg_5_9 <= _T_22578[9];
    conflictPReg_5_10 <= _T_22578[10];
    conflictPReg_5_11 <= _T_22578[11];
    conflictPReg_5_12 <= _T_22578[12];
    conflictPReg_5_13 <= _T_22578[13];
    conflictPReg_5_14 <= _T_22578[14];
    conflictPReg_5_15 <= _T_22578[15];
    conflictPReg_6_0 <= _T_23436[0];
    conflictPReg_6_1 <= _T_23436[1];
    conflictPReg_6_2 <= _T_23436[2];
    conflictPReg_6_3 <= _T_23436[3];
    conflictPReg_6_4 <= _T_23436[4];
    conflictPReg_6_5 <= _T_23436[5];
    conflictPReg_6_6 <= _T_23436[6];
    conflictPReg_6_7 <= _T_23436[7];
    conflictPReg_6_8 <= _T_23436[8];
    conflictPReg_6_9 <= _T_23436[9];
    conflictPReg_6_10 <= _T_23436[10];
    conflictPReg_6_11 <= _T_23436[11];
    conflictPReg_6_12 <= _T_23436[12];
    conflictPReg_6_13 <= _T_23436[13];
    conflictPReg_6_14 <= _T_23436[14];
    conflictPReg_6_15 <= _T_23436[15];
    conflictPReg_7_0 <= _T_24294[0];
    conflictPReg_7_1 <= _T_24294[1];
    conflictPReg_7_2 <= _T_24294[2];
    conflictPReg_7_3 <= _T_24294[3];
    conflictPReg_7_4 <= _T_24294[4];
    conflictPReg_7_5 <= _T_24294[5];
    conflictPReg_7_6 <= _T_24294[6];
    conflictPReg_7_7 <= _T_24294[7];
    conflictPReg_7_8 <= _T_24294[8];
    conflictPReg_7_9 <= _T_24294[9];
    conflictPReg_7_10 <= _T_24294[10];
    conflictPReg_7_11 <= _T_24294[11];
    conflictPReg_7_12 <= _T_24294[12];
    conflictPReg_7_13 <= _T_24294[13];
    conflictPReg_7_14 <= _T_24294[14];
    conflictPReg_7_15 <= _T_24294[15];
    conflictPReg_8_0 <= _T_25152[0];
    conflictPReg_8_1 <= _T_25152[1];
    conflictPReg_8_2 <= _T_25152[2];
    conflictPReg_8_3 <= _T_25152[3];
    conflictPReg_8_4 <= _T_25152[4];
    conflictPReg_8_5 <= _T_25152[5];
    conflictPReg_8_6 <= _T_25152[6];
    conflictPReg_8_7 <= _T_25152[7];
    conflictPReg_8_8 <= _T_25152[8];
    conflictPReg_8_9 <= _T_25152[9];
    conflictPReg_8_10 <= _T_25152[10];
    conflictPReg_8_11 <= _T_25152[11];
    conflictPReg_8_12 <= _T_25152[12];
    conflictPReg_8_13 <= _T_25152[13];
    conflictPReg_8_14 <= _T_25152[14];
    conflictPReg_8_15 <= _T_25152[15];
    conflictPReg_9_0 <= _T_26010[0];
    conflictPReg_9_1 <= _T_26010[1];
    conflictPReg_9_2 <= _T_26010[2];
    conflictPReg_9_3 <= _T_26010[3];
    conflictPReg_9_4 <= _T_26010[4];
    conflictPReg_9_5 <= _T_26010[5];
    conflictPReg_9_6 <= _T_26010[6];
    conflictPReg_9_7 <= _T_26010[7];
    conflictPReg_9_8 <= _T_26010[8];
    conflictPReg_9_9 <= _T_26010[9];
    conflictPReg_9_10 <= _T_26010[10];
    conflictPReg_9_11 <= _T_26010[11];
    conflictPReg_9_12 <= _T_26010[12];
    conflictPReg_9_13 <= _T_26010[13];
    conflictPReg_9_14 <= _T_26010[14];
    conflictPReg_9_15 <= _T_26010[15];
    conflictPReg_10_0 <= _T_26868[0];
    conflictPReg_10_1 <= _T_26868[1];
    conflictPReg_10_2 <= _T_26868[2];
    conflictPReg_10_3 <= _T_26868[3];
    conflictPReg_10_4 <= _T_26868[4];
    conflictPReg_10_5 <= _T_26868[5];
    conflictPReg_10_6 <= _T_26868[6];
    conflictPReg_10_7 <= _T_26868[7];
    conflictPReg_10_8 <= _T_26868[8];
    conflictPReg_10_9 <= _T_26868[9];
    conflictPReg_10_10 <= _T_26868[10];
    conflictPReg_10_11 <= _T_26868[11];
    conflictPReg_10_12 <= _T_26868[12];
    conflictPReg_10_13 <= _T_26868[13];
    conflictPReg_10_14 <= _T_26868[14];
    conflictPReg_10_15 <= _T_26868[15];
    conflictPReg_11_0 <= _T_27726[0];
    conflictPReg_11_1 <= _T_27726[1];
    conflictPReg_11_2 <= _T_27726[2];
    conflictPReg_11_3 <= _T_27726[3];
    conflictPReg_11_4 <= _T_27726[4];
    conflictPReg_11_5 <= _T_27726[5];
    conflictPReg_11_6 <= _T_27726[6];
    conflictPReg_11_7 <= _T_27726[7];
    conflictPReg_11_8 <= _T_27726[8];
    conflictPReg_11_9 <= _T_27726[9];
    conflictPReg_11_10 <= _T_27726[10];
    conflictPReg_11_11 <= _T_27726[11];
    conflictPReg_11_12 <= _T_27726[12];
    conflictPReg_11_13 <= _T_27726[13];
    conflictPReg_11_14 <= _T_27726[14];
    conflictPReg_11_15 <= _T_27726[15];
    conflictPReg_12_0 <= _T_28584[0];
    conflictPReg_12_1 <= _T_28584[1];
    conflictPReg_12_2 <= _T_28584[2];
    conflictPReg_12_3 <= _T_28584[3];
    conflictPReg_12_4 <= _T_28584[4];
    conflictPReg_12_5 <= _T_28584[5];
    conflictPReg_12_6 <= _T_28584[6];
    conflictPReg_12_7 <= _T_28584[7];
    conflictPReg_12_8 <= _T_28584[8];
    conflictPReg_12_9 <= _T_28584[9];
    conflictPReg_12_10 <= _T_28584[10];
    conflictPReg_12_11 <= _T_28584[11];
    conflictPReg_12_12 <= _T_28584[12];
    conflictPReg_12_13 <= _T_28584[13];
    conflictPReg_12_14 <= _T_28584[14];
    conflictPReg_12_15 <= _T_28584[15];
    conflictPReg_13_0 <= _T_29442[0];
    conflictPReg_13_1 <= _T_29442[1];
    conflictPReg_13_2 <= _T_29442[2];
    conflictPReg_13_3 <= _T_29442[3];
    conflictPReg_13_4 <= _T_29442[4];
    conflictPReg_13_5 <= _T_29442[5];
    conflictPReg_13_6 <= _T_29442[6];
    conflictPReg_13_7 <= _T_29442[7];
    conflictPReg_13_8 <= _T_29442[8];
    conflictPReg_13_9 <= _T_29442[9];
    conflictPReg_13_10 <= _T_29442[10];
    conflictPReg_13_11 <= _T_29442[11];
    conflictPReg_13_12 <= _T_29442[12];
    conflictPReg_13_13 <= _T_29442[13];
    conflictPReg_13_14 <= _T_29442[14];
    conflictPReg_13_15 <= _T_29442[15];
    conflictPReg_14_0 <= _T_30300[0];
    conflictPReg_14_1 <= _T_30300[1];
    conflictPReg_14_2 <= _T_30300[2];
    conflictPReg_14_3 <= _T_30300[3];
    conflictPReg_14_4 <= _T_30300[4];
    conflictPReg_14_5 <= _T_30300[5];
    conflictPReg_14_6 <= _T_30300[6];
    conflictPReg_14_7 <= _T_30300[7];
    conflictPReg_14_8 <= _T_30300[8];
    conflictPReg_14_9 <= _T_30300[9];
    conflictPReg_14_10 <= _T_30300[10];
    conflictPReg_14_11 <= _T_30300[11];
    conflictPReg_14_12 <= _T_30300[12];
    conflictPReg_14_13 <= _T_30300[13];
    conflictPReg_14_14 <= _T_30300[14];
    conflictPReg_14_15 <= _T_30300[15];
    conflictPReg_15_0 <= _T_31158[0];
    conflictPReg_15_1 <= _T_31158[1];
    conflictPReg_15_2 <= _T_31158[2];
    conflictPReg_15_3 <= _T_31158[3];
    conflictPReg_15_4 <= _T_31158[4];
    conflictPReg_15_5 <= _T_31158[5];
    conflictPReg_15_6 <= _T_31158[6];
    conflictPReg_15_7 <= _T_31158[7];
    conflictPReg_15_8 <= _T_31158[8];
    conflictPReg_15_9 <= _T_31158[9];
    conflictPReg_15_10 <= _T_31158[10];
    conflictPReg_15_11 <= _T_31158[11];
    conflictPReg_15_12 <= _T_31158[12];
    conflictPReg_15_13 <= _T_31158[13];
    conflictPReg_15_14 <= _T_31158[14];
    conflictPReg_15_15 <= _T_31158[15];
    storeAddrNotKnownFlagsPReg_0_0 <= _T_52612[0];
    storeAddrNotKnownFlagsPReg_0_1 <= _T_52612[1];
    storeAddrNotKnownFlagsPReg_0_2 <= _T_52612[2];
    storeAddrNotKnownFlagsPReg_0_3 <= _T_52612[3];
    storeAddrNotKnownFlagsPReg_0_4 <= _T_52612[4];
    storeAddrNotKnownFlagsPReg_0_5 <= _T_52612[5];
    storeAddrNotKnownFlagsPReg_0_6 <= _T_52612[6];
    storeAddrNotKnownFlagsPReg_0_7 <= _T_52612[7];
    storeAddrNotKnownFlagsPReg_0_8 <= _T_52612[8];
    storeAddrNotKnownFlagsPReg_0_9 <= _T_52612[9];
    storeAddrNotKnownFlagsPReg_0_10 <= _T_52612[10];
    storeAddrNotKnownFlagsPReg_0_11 <= _T_52612[11];
    storeAddrNotKnownFlagsPReg_0_12 <= _T_52612[12];
    storeAddrNotKnownFlagsPReg_0_13 <= _T_52612[13];
    storeAddrNotKnownFlagsPReg_0_14 <= _T_52612[14];
    storeAddrNotKnownFlagsPReg_0_15 <= _T_52612[15];
    storeAddrNotKnownFlagsPReg_1_0 <= _T_53470[0];
    storeAddrNotKnownFlagsPReg_1_1 <= _T_53470[1];
    storeAddrNotKnownFlagsPReg_1_2 <= _T_53470[2];
    storeAddrNotKnownFlagsPReg_1_3 <= _T_53470[3];
    storeAddrNotKnownFlagsPReg_1_4 <= _T_53470[4];
    storeAddrNotKnownFlagsPReg_1_5 <= _T_53470[5];
    storeAddrNotKnownFlagsPReg_1_6 <= _T_53470[6];
    storeAddrNotKnownFlagsPReg_1_7 <= _T_53470[7];
    storeAddrNotKnownFlagsPReg_1_8 <= _T_53470[8];
    storeAddrNotKnownFlagsPReg_1_9 <= _T_53470[9];
    storeAddrNotKnownFlagsPReg_1_10 <= _T_53470[10];
    storeAddrNotKnownFlagsPReg_1_11 <= _T_53470[11];
    storeAddrNotKnownFlagsPReg_1_12 <= _T_53470[12];
    storeAddrNotKnownFlagsPReg_1_13 <= _T_53470[13];
    storeAddrNotKnownFlagsPReg_1_14 <= _T_53470[14];
    storeAddrNotKnownFlagsPReg_1_15 <= _T_53470[15];
    storeAddrNotKnownFlagsPReg_2_0 <= _T_54328[0];
    storeAddrNotKnownFlagsPReg_2_1 <= _T_54328[1];
    storeAddrNotKnownFlagsPReg_2_2 <= _T_54328[2];
    storeAddrNotKnownFlagsPReg_2_3 <= _T_54328[3];
    storeAddrNotKnownFlagsPReg_2_4 <= _T_54328[4];
    storeAddrNotKnownFlagsPReg_2_5 <= _T_54328[5];
    storeAddrNotKnownFlagsPReg_2_6 <= _T_54328[6];
    storeAddrNotKnownFlagsPReg_2_7 <= _T_54328[7];
    storeAddrNotKnownFlagsPReg_2_8 <= _T_54328[8];
    storeAddrNotKnownFlagsPReg_2_9 <= _T_54328[9];
    storeAddrNotKnownFlagsPReg_2_10 <= _T_54328[10];
    storeAddrNotKnownFlagsPReg_2_11 <= _T_54328[11];
    storeAddrNotKnownFlagsPReg_2_12 <= _T_54328[12];
    storeAddrNotKnownFlagsPReg_2_13 <= _T_54328[13];
    storeAddrNotKnownFlagsPReg_2_14 <= _T_54328[14];
    storeAddrNotKnownFlagsPReg_2_15 <= _T_54328[15];
    storeAddrNotKnownFlagsPReg_3_0 <= _T_55186[0];
    storeAddrNotKnownFlagsPReg_3_1 <= _T_55186[1];
    storeAddrNotKnownFlagsPReg_3_2 <= _T_55186[2];
    storeAddrNotKnownFlagsPReg_3_3 <= _T_55186[3];
    storeAddrNotKnownFlagsPReg_3_4 <= _T_55186[4];
    storeAddrNotKnownFlagsPReg_3_5 <= _T_55186[5];
    storeAddrNotKnownFlagsPReg_3_6 <= _T_55186[6];
    storeAddrNotKnownFlagsPReg_3_7 <= _T_55186[7];
    storeAddrNotKnownFlagsPReg_3_8 <= _T_55186[8];
    storeAddrNotKnownFlagsPReg_3_9 <= _T_55186[9];
    storeAddrNotKnownFlagsPReg_3_10 <= _T_55186[10];
    storeAddrNotKnownFlagsPReg_3_11 <= _T_55186[11];
    storeAddrNotKnownFlagsPReg_3_12 <= _T_55186[12];
    storeAddrNotKnownFlagsPReg_3_13 <= _T_55186[13];
    storeAddrNotKnownFlagsPReg_3_14 <= _T_55186[14];
    storeAddrNotKnownFlagsPReg_3_15 <= _T_55186[15];
    storeAddrNotKnownFlagsPReg_4_0 <= _T_56044[0];
    storeAddrNotKnownFlagsPReg_4_1 <= _T_56044[1];
    storeAddrNotKnownFlagsPReg_4_2 <= _T_56044[2];
    storeAddrNotKnownFlagsPReg_4_3 <= _T_56044[3];
    storeAddrNotKnownFlagsPReg_4_4 <= _T_56044[4];
    storeAddrNotKnownFlagsPReg_4_5 <= _T_56044[5];
    storeAddrNotKnownFlagsPReg_4_6 <= _T_56044[6];
    storeAddrNotKnownFlagsPReg_4_7 <= _T_56044[7];
    storeAddrNotKnownFlagsPReg_4_8 <= _T_56044[8];
    storeAddrNotKnownFlagsPReg_4_9 <= _T_56044[9];
    storeAddrNotKnownFlagsPReg_4_10 <= _T_56044[10];
    storeAddrNotKnownFlagsPReg_4_11 <= _T_56044[11];
    storeAddrNotKnownFlagsPReg_4_12 <= _T_56044[12];
    storeAddrNotKnownFlagsPReg_4_13 <= _T_56044[13];
    storeAddrNotKnownFlagsPReg_4_14 <= _T_56044[14];
    storeAddrNotKnownFlagsPReg_4_15 <= _T_56044[15];
    storeAddrNotKnownFlagsPReg_5_0 <= _T_56902[0];
    storeAddrNotKnownFlagsPReg_5_1 <= _T_56902[1];
    storeAddrNotKnownFlagsPReg_5_2 <= _T_56902[2];
    storeAddrNotKnownFlagsPReg_5_3 <= _T_56902[3];
    storeAddrNotKnownFlagsPReg_5_4 <= _T_56902[4];
    storeAddrNotKnownFlagsPReg_5_5 <= _T_56902[5];
    storeAddrNotKnownFlagsPReg_5_6 <= _T_56902[6];
    storeAddrNotKnownFlagsPReg_5_7 <= _T_56902[7];
    storeAddrNotKnownFlagsPReg_5_8 <= _T_56902[8];
    storeAddrNotKnownFlagsPReg_5_9 <= _T_56902[9];
    storeAddrNotKnownFlagsPReg_5_10 <= _T_56902[10];
    storeAddrNotKnownFlagsPReg_5_11 <= _T_56902[11];
    storeAddrNotKnownFlagsPReg_5_12 <= _T_56902[12];
    storeAddrNotKnownFlagsPReg_5_13 <= _T_56902[13];
    storeAddrNotKnownFlagsPReg_5_14 <= _T_56902[14];
    storeAddrNotKnownFlagsPReg_5_15 <= _T_56902[15];
    storeAddrNotKnownFlagsPReg_6_0 <= _T_57760[0];
    storeAddrNotKnownFlagsPReg_6_1 <= _T_57760[1];
    storeAddrNotKnownFlagsPReg_6_2 <= _T_57760[2];
    storeAddrNotKnownFlagsPReg_6_3 <= _T_57760[3];
    storeAddrNotKnownFlagsPReg_6_4 <= _T_57760[4];
    storeAddrNotKnownFlagsPReg_6_5 <= _T_57760[5];
    storeAddrNotKnownFlagsPReg_6_6 <= _T_57760[6];
    storeAddrNotKnownFlagsPReg_6_7 <= _T_57760[7];
    storeAddrNotKnownFlagsPReg_6_8 <= _T_57760[8];
    storeAddrNotKnownFlagsPReg_6_9 <= _T_57760[9];
    storeAddrNotKnownFlagsPReg_6_10 <= _T_57760[10];
    storeAddrNotKnownFlagsPReg_6_11 <= _T_57760[11];
    storeAddrNotKnownFlagsPReg_6_12 <= _T_57760[12];
    storeAddrNotKnownFlagsPReg_6_13 <= _T_57760[13];
    storeAddrNotKnownFlagsPReg_6_14 <= _T_57760[14];
    storeAddrNotKnownFlagsPReg_6_15 <= _T_57760[15];
    storeAddrNotKnownFlagsPReg_7_0 <= _T_58618[0];
    storeAddrNotKnownFlagsPReg_7_1 <= _T_58618[1];
    storeAddrNotKnownFlagsPReg_7_2 <= _T_58618[2];
    storeAddrNotKnownFlagsPReg_7_3 <= _T_58618[3];
    storeAddrNotKnownFlagsPReg_7_4 <= _T_58618[4];
    storeAddrNotKnownFlagsPReg_7_5 <= _T_58618[5];
    storeAddrNotKnownFlagsPReg_7_6 <= _T_58618[6];
    storeAddrNotKnownFlagsPReg_7_7 <= _T_58618[7];
    storeAddrNotKnownFlagsPReg_7_8 <= _T_58618[8];
    storeAddrNotKnownFlagsPReg_7_9 <= _T_58618[9];
    storeAddrNotKnownFlagsPReg_7_10 <= _T_58618[10];
    storeAddrNotKnownFlagsPReg_7_11 <= _T_58618[11];
    storeAddrNotKnownFlagsPReg_7_12 <= _T_58618[12];
    storeAddrNotKnownFlagsPReg_7_13 <= _T_58618[13];
    storeAddrNotKnownFlagsPReg_7_14 <= _T_58618[14];
    storeAddrNotKnownFlagsPReg_7_15 <= _T_58618[15];
    storeAddrNotKnownFlagsPReg_8_0 <= _T_59476[0];
    storeAddrNotKnownFlagsPReg_8_1 <= _T_59476[1];
    storeAddrNotKnownFlagsPReg_8_2 <= _T_59476[2];
    storeAddrNotKnownFlagsPReg_8_3 <= _T_59476[3];
    storeAddrNotKnownFlagsPReg_8_4 <= _T_59476[4];
    storeAddrNotKnownFlagsPReg_8_5 <= _T_59476[5];
    storeAddrNotKnownFlagsPReg_8_6 <= _T_59476[6];
    storeAddrNotKnownFlagsPReg_8_7 <= _T_59476[7];
    storeAddrNotKnownFlagsPReg_8_8 <= _T_59476[8];
    storeAddrNotKnownFlagsPReg_8_9 <= _T_59476[9];
    storeAddrNotKnownFlagsPReg_8_10 <= _T_59476[10];
    storeAddrNotKnownFlagsPReg_8_11 <= _T_59476[11];
    storeAddrNotKnownFlagsPReg_8_12 <= _T_59476[12];
    storeAddrNotKnownFlagsPReg_8_13 <= _T_59476[13];
    storeAddrNotKnownFlagsPReg_8_14 <= _T_59476[14];
    storeAddrNotKnownFlagsPReg_8_15 <= _T_59476[15];
    storeAddrNotKnownFlagsPReg_9_0 <= _T_60334[0];
    storeAddrNotKnownFlagsPReg_9_1 <= _T_60334[1];
    storeAddrNotKnownFlagsPReg_9_2 <= _T_60334[2];
    storeAddrNotKnownFlagsPReg_9_3 <= _T_60334[3];
    storeAddrNotKnownFlagsPReg_9_4 <= _T_60334[4];
    storeAddrNotKnownFlagsPReg_9_5 <= _T_60334[5];
    storeAddrNotKnownFlagsPReg_9_6 <= _T_60334[6];
    storeAddrNotKnownFlagsPReg_9_7 <= _T_60334[7];
    storeAddrNotKnownFlagsPReg_9_8 <= _T_60334[8];
    storeAddrNotKnownFlagsPReg_9_9 <= _T_60334[9];
    storeAddrNotKnownFlagsPReg_9_10 <= _T_60334[10];
    storeAddrNotKnownFlagsPReg_9_11 <= _T_60334[11];
    storeAddrNotKnownFlagsPReg_9_12 <= _T_60334[12];
    storeAddrNotKnownFlagsPReg_9_13 <= _T_60334[13];
    storeAddrNotKnownFlagsPReg_9_14 <= _T_60334[14];
    storeAddrNotKnownFlagsPReg_9_15 <= _T_60334[15];
    storeAddrNotKnownFlagsPReg_10_0 <= _T_61192[0];
    storeAddrNotKnownFlagsPReg_10_1 <= _T_61192[1];
    storeAddrNotKnownFlagsPReg_10_2 <= _T_61192[2];
    storeAddrNotKnownFlagsPReg_10_3 <= _T_61192[3];
    storeAddrNotKnownFlagsPReg_10_4 <= _T_61192[4];
    storeAddrNotKnownFlagsPReg_10_5 <= _T_61192[5];
    storeAddrNotKnownFlagsPReg_10_6 <= _T_61192[6];
    storeAddrNotKnownFlagsPReg_10_7 <= _T_61192[7];
    storeAddrNotKnownFlagsPReg_10_8 <= _T_61192[8];
    storeAddrNotKnownFlagsPReg_10_9 <= _T_61192[9];
    storeAddrNotKnownFlagsPReg_10_10 <= _T_61192[10];
    storeAddrNotKnownFlagsPReg_10_11 <= _T_61192[11];
    storeAddrNotKnownFlagsPReg_10_12 <= _T_61192[12];
    storeAddrNotKnownFlagsPReg_10_13 <= _T_61192[13];
    storeAddrNotKnownFlagsPReg_10_14 <= _T_61192[14];
    storeAddrNotKnownFlagsPReg_10_15 <= _T_61192[15];
    storeAddrNotKnownFlagsPReg_11_0 <= _T_62050[0];
    storeAddrNotKnownFlagsPReg_11_1 <= _T_62050[1];
    storeAddrNotKnownFlagsPReg_11_2 <= _T_62050[2];
    storeAddrNotKnownFlagsPReg_11_3 <= _T_62050[3];
    storeAddrNotKnownFlagsPReg_11_4 <= _T_62050[4];
    storeAddrNotKnownFlagsPReg_11_5 <= _T_62050[5];
    storeAddrNotKnownFlagsPReg_11_6 <= _T_62050[6];
    storeAddrNotKnownFlagsPReg_11_7 <= _T_62050[7];
    storeAddrNotKnownFlagsPReg_11_8 <= _T_62050[8];
    storeAddrNotKnownFlagsPReg_11_9 <= _T_62050[9];
    storeAddrNotKnownFlagsPReg_11_10 <= _T_62050[10];
    storeAddrNotKnownFlagsPReg_11_11 <= _T_62050[11];
    storeAddrNotKnownFlagsPReg_11_12 <= _T_62050[12];
    storeAddrNotKnownFlagsPReg_11_13 <= _T_62050[13];
    storeAddrNotKnownFlagsPReg_11_14 <= _T_62050[14];
    storeAddrNotKnownFlagsPReg_11_15 <= _T_62050[15];
    storeAddrNotKnownFlagsPReg_12_0 <= _T_62908[0];
    storeAddrNotKnownFlagsPReg_12_1 <= _T_62908[1];
    storeAddrNotKnownFlagsPReg_12_2 <= _T_62908[2];
    storeAddrNotKnownFlagsPReg_12_3 <= _T_62908[3];
    storeAddrNotKnownFlagsPReg_12_4 <= _T_62908[4];
    storeAddrNotKnownFlagsPReg_12_5 <= _T_62908[5];
    storeAddrNotKnownFlagsPReg_12_6 <= _T_62908[6];
    storeAddrNotKnownFlagsPReg_12_7 <= _T_62908[7];
    storeAddrNotKnownFlagsPReg_12_8 <= _T_62908[8];
    storeAddrNotKnownFlagsPReg_12_9 <= _T_62908[9];
    storeAddrNotKnownFlagsPReg_12_10 <= _T_62908[10];
    storeAddrNotKnownFlagsPReg_12_11 <= _T_62908[11];
    storeAddrNotKnownFlagsPReg_12_12 <= _T_62908[12];
    storeAddrNotKnownFlagsPReg_12_13 <= _T_62908[13];
    storeAddrNotKnownFlagsPReg_12_14 <= _T_62908[14];
    storeAddrNotKnownFlagsPReg_12_15 <= _T_62908[15];
    storeAddrNotKnownFlagsPReg_13_0 <= _T_63766[0];
    storeAddrNotKnownFlagsPReg_13_1 <= _T_63766[1];
    storeAddrNotKnownFlagsPReg_13_2 <= _T_63766[2];
    storeAddrNotKnownFlagsPReg_13_3 <= _T_63766[3];
    storeAddrNotKnownFlagsPReg_13_4 <= _T_63766[4];
    storeAddrNotKnownFlagsPReg_13_5 <= _T_63766[5];
    storeAddrNotKnownFlagsPReg_13_6 <= _T_63766[6];
    storeAddrNotKnownFlagsPReg_13_7 <= _T_63766[7];
    storeAddrNotKnownFlagsPReg_13_8 <= _T_63766[8];
    storeAddrNotKnownFlagsPReg_13_9 <= _T_63766[9];
    storeAddrNotKnownFlagsPReg_13_10 <= _T_63766[10];
    storeAddrNotKnownFlagsPReg_13_11 <= _T_63766[11];
    storeAddrNotKnownFlagsPReg_13_12 <= _T_63766[12];
    storeAddrNotKnownFlagsPReg_13_13 <= _T_63766[13];
    storeAddrNotKnownFlagsPReg_13_14 <= _T_63766[14];
    storeAddrNotKnownFlagsPReg_13_15 <= _T_63766[15];
    storeAddrNotKnownFlagsPReg_14_0 <= _T_64624[0];
    storeAddrNotKnownFlagsPReg_14_1 <= _T_64624[1];
    storeAddrNotKnownFlagsPReg_14_2 <= _T_64624[2];
    storeAddrNotKnownFlagsPReg_14_3 <= _T_64624[3];
    storeAddrNotKnownFlagsPReg_14_4 <= _T_64624[4];
    storeAddrNotKnownFlagsPReg_14_5 <= _T_64624[5];
    storeAddrNotKnownFlagsPReg_14_6 <= _T_64624[6];
    storeAddrNotKnownFlagsPReg_14_7 <= _T_64624[7];
    storeAddrNotKnownFlagsPReg_14_8 <= _T_64624[8];
    storeAddrNotKnownFlagsPReg_14_9 <= _T_64624[9];
    storeAddrNotKnownFlagsPReg_14_10 <= _T_64624[10];
    storeAddrNotKnownFlagsPReg_14_11 <= _T_64624[11];
    storeAddrNotKnownFlagsPReg_14_12 <= _T_64624[12];
    storeAddrNotKnownFlagsPReg_14_13 <= _T_64624[13];
    storeAddrNotKnownFlagsPReg_14_14 <= _T_64624[14];
    storeAddrNotKnownFlagsPReg_14_15 <= _T_64624[15];
    storeAddrNotKnownFlagsPReg_15_0 <= _T_65482[0];
    storeAddrNotKnownFlagsPReg_15_1 <= _T_65482[1];
    storeAddrNotKnownFlagsPReg_15_2 <= _T_65482[2];
    storeAddrNotKnownFlagsPReg_15_3 <= _T_65482[3];
    storeAddrNotKnownFlagsPReg_15_4 <= _T_65482[4];
    storeAddrNotKnownFlagsPReg_15_5 <= _T_65482[5];
    storeAddrNotKnownFlagsPReg_15_6 <= _T_65482[6];
    storeAddrNotKnownFlagsPReg_15_7 <= _T_65482[7];
    storeAddrNotKnownFlagsPReg_15_8 <= _T_65482[8];
    storeAddrNotKnownFlagsPReg_15_9 <= _T_65482[9];
    storeAddrNotKnownFlagsPReg_15_10 <= _T_65482[10];
    storeAddrNotKnownFlagsPReg_15_11 <= _T_65482[11];
    storeAddrNotKnownFlagsPReg_15_12 <= _T_65482[12];
    storeAddrNotKnownFlagsPReg_15_13 <= _T_65482[13];
    storeAddrNotKnownFlagsPReg_15_14 <= _T_65482[14];
    storeAddrNotKnownFlagsPReg_15_15 <= _T_65482[15];
    shiftedStoreDataKnownPReg_0 <= _T_5978[0];
    shiftedStoreDataKnownPReg_1 <= _T_5978[1];
    shiftedStoreDataKnownPReg_2 <= _T_5978[2];
    shiftedStoreDataKnownPReg_3 <= _T_5978[3];
    shiftedStoreDataKnownPReg_4 <= _T_5978[4];
    shiftedStoreDataKnownPReg_5 <= _T_5978[5];
    shiftedStoreDataKnownPReg_6 <= _T_5978[6];
    shiftedStoreDataKnownPReg_7 <= _T_5978[7];
    shiftedStoreDataKnownPReg_8 <= _T_5978[8];
    shiftedStoreDataKnownPReg_9 <= _T_5978[9];
    shiftedStoreDataKnownPReg_10 <= _T_5978[10];
    shiftedStoreDataKnownPReg_11 <= _T_5978[11];
    shiftedStoreDataKnownPReg_12 <= _T_5978[12];
    shiftedStoreDataKnownPReg_13 <= _T_5978[13];
    shiftedStoreDataKnownPReg_14 <= _T_5978[14];
    shiftedStoreDataKnownPReg_15 <= _T_5978[15];
    shiftedStoreDataQPreg_0 <= _T_5121[31:0];
    shiftedStoreDataQPreg_1 <= _T_5121[63:32];
    shiftedStoreDataQPreg_2 <= _T_5121[95:64];
    shiftedStoreDataQPreg_3 <= _T_5121[127:96];
    shiftedStoreDataQPreg_4 <= _T_5121[159:128];
    shiftedStoreDataQPreg_5 <= _T_5121[191:160];
    shiftedStoreDataQPreg_6 <= _T_5121[223:192];
    shiftedStoreDataQPreg_7 <= _T_5121[255:224];
    shiftedStoreDataQPreg_8 <= _T_5121[287:256];
    shiftedStoreDataQPreg_9 <= _T_5121[319:288];
    shiftedStoreDataQPreg_10 <= _T_5121[351:320];
    shiftedStoreDataQPreg_11 <= _T_5121[383:352];
    shiftedStoreDataQPreg_12 <= _T_5121[415:384];
    shiftedStoreDataQPreg_13 <= _T_5121[447:416];
    shiftedStoreDataQPreg_14 <= _T_5121[479:448];
    shiftedStoreDataQPreg_15 <= _T_5121[511:480];
    addrKnownPReg_0 <= addrKnown_0;
    addrKnownPReg_1 <= addrKnown_1;
    addrKnownPReg_2 <= addrKnown_2;
    addrKnownPReg_3 <= addrKnown_3;
    addrKnownPReg_4 <= addrKnown_4;
    addrKnownPReg_5 <= addrKnown_5;
    addrKnownPReg_6 <= addrKnown_6;
    addrKnownPReg_7 <= addrKnown_7;
    addrKnownPReg_8 <= addrKnown_8;
    addrKnownPReg_9 <= addrKnown_9;
    addrKnownPReg_10 <= addrKnown_10;
    addrKnownPReg_11 <= addrKnown_11;
    addrKnownPReg_12 <= addrKnown_12;
    addrKnownPReg_13 <= addrKnown_13;
    addrKnownPReg_14 <= addrKnown_14;
    addrKnownPReg_15 <= addrKnown_15;
    dataKnownPReg_0 <= dataKnown_0;
    dataKnownPReg_1 <= dataKnown_1;
    dataKnownPReg_2 <= dataKnown_2;
    dataKnownPReg_3 <= dataKnown_3;
    dataKnownPReg_4 <= dataKnown_4;
    dataKnownPReg_5 <= dataKnown_5;
    dataKnownPReg_6 <= dataKnown_6;
    dataKnownPReg_7 <= dataKnown_7;
    dataKnownPReg_8 <= dataKnown_8;
    dataKnownPReg_9 <= dataKnown_9;
    dataKnownPReg_10 <= dataKnown_10;
    dataKnownPReg_11 <= dataKnown_11;
    dataKnownPReg_12 <= dataKnown_12;
    dataKnownPReg_13 <= dataKnown_13;
    dataKnownPReg_14 <= dataKnown_14;
    dataKnownPReg_15 <= dataKnown_15;
    if (reset) begin
      loadInitiated_15 <= 1'h0;
    end else begin
      if (initBits_15) begin
        loadInitiated_15 <= 1'h0;
      end else begin
        if (_T_92231) begin
          loadInitiated_15 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_14 <= 1'h0;
    end else begin
      if (initBits_14) begin
        loadInitiated_14 <= 1'h0;
      end else begin
        if (_T_92228) begin
          loadInitiated_14 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_13 <= 1'h0;
    end else begin
      if (initBits_13) begin
        loadInitiated_13 <= 1'h0;
      end else begin
        if (_T_92225) begin
          loadInitiated_13 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_12 <= 1'h0;
    end else begin
      if (initBits_12) begin
        loadInitiated_12 <= 1'h0;
      end else begin
        if (_T_92222) begin
          loadInitiated_12 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_11 <= 1'h0;
    end else begin
      if (initBits_11) begin
        loadInitiated_11 <= 1'h0;
      end else begin
        if (_T_92219) begin
          loadInitiated_11 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_10 <= 1'h0;
    end else begin
      if (initBits_10) begin
        loadInitiated_10 <= 1'h0;
      end else begin
        if (_T_92216) begin
          loadInitiated_10 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_9 <= 1'h0;
    end else begin
      if (initBits_9) begin
        loadInitiated_9 <= 1'h0;
      end else begin
        if (_T_92213) begin
          loadInitiated_9 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_8 <= 1'h0;
    end else begin
      if (initBits_8) begin
        loadInitiated_8 <= 1'h0;
      end else begin
        if (_T_92210) begin
          loadInitiated_8 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_7 <= 1'h0;
    end else begin
      if (initBits_7) begin
        loadInitiated_7 <= 1'h0;
      end else begin
        if (_T_92207) begin
          loadInitiated_7 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_6 <= 1'h0;
    end else begin
      if (initBits_6) begin
        loadInitiated_6 <= 1'h0;
      end else begin
        if (_T_92204) begin
          loadInitiated_6 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_5 <= 1'h0;
    end else begin
      if (initBits_5) begin
        loadInitiated_5 <= 1'h0;
      end else begin
        if (_T_92201) begin
          loadInitiated_5 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_4 <= 1'h0;
    end else begin
      if (initBits_4) begin
        loadInitiated_4 <= 1'h0;
      end else begin
        if (_T_92198) begin
          loadInitiated_4 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_3 <= 1'h0;
    end else begin
      if (initBits_3) begin
        loadInitiated_3 <= 1'h0;
      end else begin
        if (_T_92195) begin
          loadInitiated_3 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_2 <= 1'h0;
    end else begin
      if (initBits_2) begin
        loadInitiated_2 <= 1'h0;
      end else begin
        if (_T_92192) begin
          loadInitiated_2 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_1 <= 1'h0;
    end else begin
      if (initBits_1) begin
        loadInitiated_1 <= 1'h0;
      end else begin
        if (_T_92189) begin
          loadInitiated_1 <= 1'h1;
        end
      end
    end
    if (reset) begin
      loadInitiated_0 <= 1'h0;
    end else begin
      if (initBits_0) begin
        loadInitiated_0 <= 1'h0;
      end else begin
        if (_T_92186) begin
          loadInitiated_0 <= 1'h1;
        end
      end
    end
  end
endmodule
module GROUP_ALLOCATOR_LSQ_a( // @[:@42581.2]
  output [3:0] io_bbLoadOffsets_0, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_1, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_2, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_3, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_4, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_5, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_6, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_7, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_8, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_9, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_10, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_11, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_12, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_13, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_14, // @[:@42584.4]
  output [3:0] io_bbLoadOffsets_15, // @[:@42584.4]
  output       io_bbNumLoads, // @[:@42584.4]
  input  [3:0] io_loadTail, // @[:@42584.4]
  input  [3:0] io_loadHead, // @[:@42584.4]
  input        io_loadEmpty, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_0, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_1, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_2, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_3, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_4, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_5, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_6, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_7, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_8, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_9, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_10, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_11, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_12, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_13, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_14, // @[:@42584.4]
  output [3:0] io_bbStoreOffsets_15, // @[:@42584.4]
  output       io_bbNumStores, // @[:@42584.4]
  input  [3:0] io_storeTail, // @[:@42584.4]
  input  [3:0] io_storeHead, // @[:@42584.4]
  input        io_storeEmpty, // @[:@42584.4]
  output       io_bbStart, // @[:@42584.4]
  input        io_bbStartSignals_0, // @[:@42584.4]
  input        io_bbStartSignals_1, // @[:@42584.4]
  output       io_readyToPrevious_0, // @[:@42584.4]
  output       io_readyToPrevious_1, // @[:@42584.4]
  output       io_loadPortsEnable_0, // @[:@42584.4]
  output       io_storePortsEnable_0 // @[:@42584.4]
);
  wire  _T_244; // @[GroupAllocator.scala 42:25:@42587.4]
  wire  _T_245; // @[GroupAllocator.scala 42:16:@42588.4]
  wire [4:0] _GEN_68; // @[GroupAllocator.scala 43:36:@42590.6]
  wire [5:0] _T_247; // @[GroupAllocator.scala 43:36:@42590.6]
  wire [5:0] _T_248; // @[GroupAllocator.scala 43:36:@42591.6]
  wire [4:0] _T_249; // @[GroupAllocator.scala 43:36:@42592.6]
  wire [4:0] _GEN_69; // @[GroupAllocator.scala 43:43:@42593.6]
  wire [5:0] _T_250; // @[GroupAllocator.scala 43:43:@42593.6]
  wire [4:0] _T_251; // @[GroupAllocator.scala 43:43:@42594.6]
  wire [4:0] _T_252; // @[GroupAllocator.scala 45:22:@42598.6]
  wire [4:0] _T_253; // @[GroupAllocator.scala 45:22:@42599.6]
  wire [3:0] _T_254; // @[GroupAllocator.scala 45:22:@42600.6]
  wire [4:0] emptyLoadSlots; // @[GroupAllocator.scala 42:34:@42589.4]
  wire  _T_256; // @[GroupAllocator.scala 42:25:@42604.4]
  wire  _T_257; // @[GroupAllocator.scala 42:16:@42605.4]
  wire [4:0] _GEN_70; // @[GroupAllocator.scala 43:36:@42607.6]
  wire [5:0] _T_259; // @[GroupAllocator.scala 43:36:@42607.6]
  wire [5:0] _T_260; // @[GroupAllocator.scala 43:36:@42608.6]
  wire [4:0] _T_261; // @[GroupAllocator.scala 43:36:@42609.6]
  wire [4:0] _GEN_71; // @[GroupAllocator.scala 43:43:@42610.6]
  wire [5:0] _T_262; // @[GroupAllocator.scala 43:43:@42610.6]
  wire [4:0] _T_263; // @[GroupAllocator.scala 43:43:@42611.6]
  wire [4:0] _T_264; // @[GroupAllocator.scala 45:22:@42615.6]
  wire [4:0] _T_265; // @[GroupAllocator.scala 45:22:@42616.6]
  wire [3:0] _T_266; // @[GroupAllocator.scala 45:22:@42617.6]
  wire [4:0] emptyStoreSlots; // @[GroupAllocator.scala 42:34:@42606.4]
  wire  possibleAllocations_0; // @[GroupAllocator.scala 56:106:@42631.4]
  wire  possibleAllocations_1; // @[GroupAllocator.scala 56:106:@42632.4]
  wire  allocatedBBIdx; // @[Mux.scala 31:69:@42636.4]
  wire  _T_300; // @[GroupAllocator.scala 69:43:@42640.4]
  wire  _T_476; // @[Mux.scala 46:16:@42789.6]
  wire [5:0] _T_898; // @[GroupAllocator.scala 110:34:@42950.6]
  wire [4:0] _T_899; // @[GroupAllocator.scala 110:34:@42951.6]
  wire [5:0] _T_901; // @[GroupAllocator.scala 110:55:@42952.6]
  wire [5:0] _T_902; // @[GroupAllocator.scala 110:55:@42953.6]
  wire [4:0] _T_903; // @[GroupAllocator.scala 110:55:@42954.6]
  wire [5:0] _T_905; // @[util.scala 10:8:@42955.6]
  wire [5:0] _GEN_0; // @[util.scala 10:14:@42956.6]
  wire [4:0] _T_906; // @[util.scala 10:14:@42956.6]
  wire [3:0] _T_1156; // @[GroupAllocator.scala 110:90:@43118.6 GroupAllocator.scala 110:90:@43119.6]
  wire [3:0] _T_1390_0; // @[Mux.scala 46:16:@43273.6]
  wire [3:0] _T_1427_0; // @[Mux.scala 46:16:@43275.6]
  wire [5:0] _T_1504; // @[GroupAllocator.scala 115:33:@43309.6]
  wire [4:0] _T_1505; // @[GroupAllocator.scala 115:33:@43310.6]
  wire [5:0] _T_1507; // @[GroupAllocator.scala 115:54:@43311.6]
  wire [5:0] _T_1508; // @[GroupAllocator.scala 115:54:@43312.6]
  wire [4:0] _T_1509; // @[GroupAllocator.scala 115:54:@43313.6]
  wire [5:0] _T_1511; // @[util.scala 10:8:@43314.6]
  wire [5:0] _GEN_1; // @[util.scala 10:14:@43315.6]
  wire [4:0] _T_1512; // @[util.scala 10:14:@43315.6]
  wire [3:0] _T_1762; // @[GroupAllocator.scala 115:89:@43477.6 GroupAllocator.scala 115:89:@43478.6]
  wire [3:0] _T_1996_0; // @[Mux.scala 46:16:@43632.6]
  wire [3:0] _T_2033_0; // @[Mux.scala 46:16:@43634.6]
  assign _T_244 = io_loadHead < io_loadTail; // @[GroupAllocator.scala 42:25:@42587.4]
  assign _T_245 = io_loadEmpty | _T_244; // @[GroupAllocator.scala 42:16:@42588.4]
  assign _GEN_68 = {{1'd0}, io_loadTail}; // @[GroupAllocator.scala 43:36:@42590.6]
  assign _T_247 = 5'h10 - _GEN_68; // @[GroupAllocator.scala 43:36:@42590.6]
  assign _T_248 = $unsigned(_T_247); // @[GroupAllocator.scala 43:36:@42591.6]
  assign _T_249 = _T_248[4:0]; // @[GroupAllocator.scala 43:36:@42592.6]
  assign _GEN_69 = {{1'd0}, io_loadHead}; // @[GroupAllocator.scala 43:43:@42593.6]
  assign _T_250 = _T_249 + _GEN_69; // @[GroupAllocator.scala 43:43:@42593.6]
  assign _T_251 = _T_249 + _GEN_69; // @[GroupAllocator.scala 43:43:@42594.6]
  assign _T_252 = io_loadHead - io_loadTail; // @[GroupAllocator.scala 45:22:@42598.6]
  assign _T_253 = $unsigned(_T_252); // @[GroupAllocator.scala 45:22:@42599.6]
  assign _T_254 = _T_253[3:0]; // @[GroupAllocator.scala 45:22:@42600.6]
  assign emptyLoadSlots = _T_245 ? _T_251 : {{1'd0}, _T_254}; // @[GroupAllocator.scala 42:34:@42589.4]
  assign _T_256 = io_storeHead < io_storeTail; // @[GroupAllocator.scala 42:25:@42604.4]
  assign _T_257 = io_storeEmpty | _T_256; // @[GroupAllocator.scala 42:16:@42605.4]
  assign _GEN_70 = {{1'd0}, io_storeTail}; // @[GroupAllocator.scala 43:36:@42607.6]
  assign _T_259 = 5'h10 - _GEN_70; // @[GroupAllocator.scala 43:36:@42607.6]
  assign _T_260 = $unsigned(_T_259); // @[GroupAllocator.scala 43:36:@42608.6]
  assign _T_261 = _T_260[4:0]; // @[GroupAllocator.scala 43:36:@42609.6]
  assign _GEN_71 = {{1'd0}, io_storeHead}; // @[GroupAllocator.scala 43:43:@42610.6]
  assign _T_262 = _T_261 + _GEN_71; // @[GroupAllocator.scala 43:43:@42610.6]
  assign _T_263 = _T_261 + _GEN_71; // @[GroupAllocator.scala 43:43:@42611.6]
  assign _T_264 = io_storeHead - io_storeTail; // @[GroupAllocator.scala 45:22:@42615.6]
  assign _T_265 = $unsigned(_T_264); // @[GroupAllocator.scala 45:22:@42616.6]
  assign _T_266 = _T_265[3:0]; // @[GroupAllocator.scala 45:22:@42617.6]
  assign emptyStoreSlots = _T_257 ? _T_263 : {{1'd0}, _T_266}; // @[GroupAllocator.scala 42:34:@42606.4]
  assign possibleAllocations_0 = io_readyToPrevious_0 & io_bbStartSignals_0; // @[GroupAllocator.scala 56:106:@42631.4]
  assign possibleAllocations_1 = io_readyToPrevious_1 & io_bbStartSignals_1; // @[GroupAllocator.scala 56:106:@42632.4]
  assign allocatedBBIdx = possibleAllocations_0 ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@42636.4]
  assign _T_300 = 1'h0 == allocatedBBIdx; // @[GroupAllocator.scala 69:43:@42640.4]
  assign _T_476 = _T_300 ? 1'h0 : allocatedBBIdx; // @[Mux.scala 46:16:@42789.6]
  assign _T_898 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@42950.6]
  assign _T_899 = _GEN_70 + 5'h10; // @[GroupAllocator.scala 110:34:@42951.6]
  assign _T_901 = _T_899 - 5'h1; // @[GroupAllocator.scala 110:55:@42952.6]
  assign _T_902 = $unsigned(_T_901); // @[GroupAllocator.scala 110:55:@42953.6]
  assign _T_903 = _T_902[4:0]; // @[GroupAllocator.scala 110:55:@42954.6]
  assign _T_905 = {{1'd0}, _T_903}; // @[util.scala 10:8:@42955.6]
  assign _GEN_0 = _T_905 % 6'h10; // @[util.scala 10:14:@42956.6]
  assign _T_906 = _GEN_0[4:0]; // @[util.scala 10:14:@42956.6]
  assign _T_1156 = _T_906[3:0]; // @[GroupAllocator.scala 110:90:@43118.6 GroupAllocator.scala 110:90:@43119.6]
  assign _T_1390_0 = allocatedBBIdx ? _T_1156 : 4'h0; // @[Mux.scala 46:16:@43273.6]
  assign _T_1427_0 = _T_300 ? _T_1156 : _T_1390_0; // @[Mux.scala 46:16:@43275.6]
  assign _T_1504 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@43309.6]
  assign _T_1505 = _GEN_68 + 5'h10; // @[GroupAllocator.scala 115:33:@43310.6]
  assign _T_1507 = _T_1505 - 5'h1; // @[GroupAllocator.scala 115:54:@43311.6]
  assign _T_1508 = $unsigned(_T_1507); // @[GroupAllocator.scala 115:54:@43312.6]
  assign _T_1509 = _T_1508[4:0]; // @[GroupAllocator.scala 115:54:@43313.6]
  assign _T_1511 = {{1'd0}, _T_1509}; // @[util.scala 10:8:@43314.6]
  assign _GEN_1 = _T_1511 % 6'h10; // @[util.scala 10:14:@43315.6]
  assign _T_1512 = _GEN_1[4:0]; // @[util.scala 10:14:@43315.6]
  assign _T_1762 = _T_1512[3:0]; // @[GroupAllocator.scala 115:89:@43477.6 GroupAllocator.scala 115:89:@43478.6]
  assign _T_1996_0 = allocatedBBIdx ? _T_1762 : 4'h0; // @[Mux.scala 46:16:@43632.6]
  assign _T_2033_0 = _T_300 ? _T_1762 : _T_1996_0; // @[Mux.scala 46:16:@43634.6]
  assign io_bbLoadOffsets_0 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42731.4 GroupAllocator.scala 106:22:@43276.6]
  assign io_bbLoadOffsets_1 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42732.4 GroupAllocator.scala 106:22:@43277.6]
  assign io_bbLoadOffsets_2 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42733.4 GroupAllocator.scala 106:22:@43278.6]
  assign io_bbLoadOffsets_3 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42734.4 GroupAllocator.scala 106:22:@43279.6]
  assign io_bbLoadOffsets_4 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42735.4 GroupAllocator.scala 106:22:@43280.6]
  assign io_bbLoadOffsets_5 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42736.4 GroupAllocator.scala 106:22:@43281.6]
  assign io_bbLoadOffsets_6 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42737.4 GroupAllocator.scala 106:22:@43282.6]
  assign io_bbLoadOffsets_7 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42738.4 GroupAllocator.scala 106:22:@43283.6]
  assign io_bbLoadOffsets_8 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42739.4 GroupAllocator.scala 106:22:@43284.6]
  assign io_bbLoadOffsets_9 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42740.4 GroupAllocator.scala 106:22:@43285.6]
  assign io_bbLoadOffsets_10 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42741.4 GroupAllocator.scala 106:22:@43286.6]
  assign io_bbLoadOffsets_11 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42742.4 GroupAllocator.scala 106:22:@43287.6]
  assign io_bbLoadOffsets_12 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42743.4 GroupAllocator.scala 106:22:@43288.6]
  assign io_bbLoadOffsets_13 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42744.4 GroupAllocator.scala 106:22:@43289.6]
  assign io_bbLoadOffsets_14 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42745.4 GroupAllocator.scala 106:22:@43290.6]
  assign io_bbLoadOffsets_15 = io_bbStart ? _T_1427_0 : 4'h0; // @[GroupAllocator.scala 89:20:@42746.4 GroupAllocator.scala 106:22:@43291.6]
  assign io_bbNumLoads = io_bbStart ? _T_300 : 1'h0; // @[GroupAllocator.scala 85:17:@42646.4 GroupAllocator.scala 93:19:@42785.6]
  assign io_bbStoreOffsets_0 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42764.4 GroupAllocator.scala 111:23:@43635.6]
  assign io_bbStoreOffsets_1 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42765.4 GroupAllocator.scala 111:23:@43636.6]
  assign io_bbStoreOffsets_2 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42766.4 GroupAllocator.scala 111:23:@43637.6]
  assign io_bbStoreOffsets_3 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42767.4 GroupAllocator.scala 111:23:@43638.6]
  assign io_bbStoreOffsets_4 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42768.4 GroupAllocator.scala 111:23:@43639.6]
  assign io_bbStoreOffsets_5 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42769.4 GroupAllocator.scala 111:23:@43640.6]
  assign io_bbStoreOffsets_6 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42770.4 GroupAllocator.scala 111:23:@43641.6]
  assign io_bbStoreOffsets_7 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42771.4 GroupAllocator.scala 111:23:@43642.6]
  assign io_bbStoreOffsets_8 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42772.4 GroupAllocator.scala 111:23:@43643.6]
  assign io_bbStoreOffsets_9 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42773.4 GroupAllocator.scala 111:23:@43644.6]
  assign io_bbStoreOffsets_10 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42774.4 GroupAllocator.scala 111:23:@43645.6]
  assign io_bbStoreOffsets_11 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42775.4 GroupAllocator.scala 111:23:@43646.6]
  assign io_bbStoreOffsets_12 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42776.4 GroupAllocator.scala 111:23:@43647.6]
  assign io_bbStoreOffsets_13 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42777.4 GroupAllocator.scala 111:23:@43648.6]
  assign io_bbStoreOffsets_14 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42778.4 GroupAllocator.scala 111:23:@43649.6]
  assign io_bbStoreOffsets_15 = io_bbStart ? _T_2033_0 : 4'h0; // @[GroupAllocator.scala 90:21:@42779.4 GroupAllocator.scala 111:23:@43650.6]
  assign io_bbNumStores = io_bbStart ? _T_476 : 1'h0; // @[GroupAllocator.scala 86:18:@42647.4 GroupAllocator.scala 94:20:@42790.6]
  assign io_bbStart = possibleAllocations_0 | possibleAllocations_1; // @[GroupAllocator.scala 59:14:@42639.4]
  assign io_readyToPrevious_0 = 5'h1 <= emptyLoadSlots; // @[GroupAllocator.scala 53:22:@42629.4]
  assign io_readyToPrevious_1 = 5'h1 <= emptyStoreSlots; // @[GroupAllocator.scala 53:22:@42630.4]
  assign io_loadPortsEnable_0 = _T_300 & io_bbStart; // @[GroupAllocator.scala 69:29:@42642.4]
  assign io_storePortsEnable_0 = allocatedBBIdx & io_bbStart; // @[GroupAllocator.scala 78:30:@42645.4]
endmodule
module AXI_WRITE( // @[:@43653.2]
  input         clock, // @[:@43654.4]
  input         reset, // @[:@43655.4]
  input  [30:0] io_storeAddrToMem, // @[:@43656.4]
  input  [31:0] io_storeDataToMem, // @[:@43656.4]
  output        io_storeQIdxInToAW_ready, // @[:@43656.4]
  input         io_storeQIdxInToAW_valid, // @[:@43656.4]
  input  [3:0]  io_storeQIdxInToAW_bits, // @[:@43656.4]
  output [3:0]  io_storeQIdxOutFromAW, // @[:@43656.4]
  output        io_storeQIdxOutFromAWValid, // @[:@43656.4]
  output        io_AWID, // @[:@43656.4]
  output [30:0] io_AWADDR, // @[:@43656.4]
  output [7:0]  io_AWLEN, // @[:@43656.4]
  output [2:0]  io_AWSIZE, // @[:@43656.4]
  output [1:0]  io_AWBURST, // @[:@43656.4]
  output [2:0]  io_AWPROT, // @[:@43656.4]
  output        io_AWVALID, // @[:@43656.4]
  input         io_AWREADY, // @[:@43656.4]
  output        io_AWLOCK, // @[:@43656.4]
  output [3:0]  io_AWCACHE, // @[:@43656.4]
  output [3:0]  io_AWQOS, // @[:@43656.4]
  output [3:0]  io_AWREGION, // @[:@43656.4]
  output        io_WID, // @[:@43656.4]
  output [31:0] io_WDATA, // @[:@43656.4]
  output [3:0]  io_WSTRB, // @[:@43656.4]
  output        io_WLAST, // @[:@43656.4]
  output        io_WVALID, // @[:@43656.4]
  input         io_WREADY, // @[:@43656.4]
  input         io_BID, // @[:@43656.4]
  input  [1:0]  io_BRESP, // @[:@43656.4]
  input         io_BVALID, // @[:@43656.4]
  output        io_BREADY // @[:@43656.4]
);
  reg [3:0] idxArray_0; // @[AxiWrite.scala 57:31:@43661.4]
  reg [31:0] _RAND_0;
  reg [3:0] idxArray_1; // @[AxiWrite.scala 57:31:@43661.4]
  reg [31:0] _RAND_1;
  reg  waitingForResponse_0; // @[AxiWrite.scala 58:41:@43665.4]
  reg [31:0] _RAND_2;
  wire  _T_126; // @[AxiWrite.scala 59:81:@43666.4]
  wire  firstFreeIdx; // @[Mux.scala 31:69:@43671.4]
  wire  _T_146; // @[AxiWrite.scala 63:62:@43676.4]
  reg [1:0] r_AW_BURST; // @[AxiWrite.scala 70:33:@43681.4]
  reg [31:0] _RAND_3;
  reg [5:0] r_AW_ADDR; // @[AxiWrite.scala 71:33:@43682.4]
  reg [31:0] _RAND_4;
  reg [7:0] r_AW_LEN; // @[AxiWrite.scala 72:33:@43683.4]
  reg [31:0] _RAND_5;
  reg [2:0] r_AW_SIZE; // @[AxiWrite.scala 73:33:@43684.4]
  reg [31:0] _RAND_6;
  reg  r_AW_ID; // @[AxiWrite.scala 74:33:@43685.4]
  reg [31:0] _RAND_7;
  reg  r_AW_VALID; // @[AxiWrite.scala 75:33:@43686.4]
  reg [31:0] _RAND_8;
  reg [2:0] r_AW_PROT; // @[AxiWrite.scala 76:33:@43687.4]
  reg [31:0] _RAND_9;
  reg [3:0] r_AW_QOS; // @[AxiWrite.scala 77:34:@43688.4]
  reg [31:0] _RAND_10;
  reg  r_AW_LOCK; // @[AxiWrite.scala 78:34:@43689.4]
  reg [31:0] _RAND_11;
  reg [3:0] r_AW_CACHE; // @[AxiWrite.scala 79:34:@43690.4]
  reg [31:0] _RAND_12;
  reg [3:0] r_AW_REGION; // @[AxiWrite.scala 80:34:@43691.4]
  reg [31:0] _RAND_13;
  reg [31:0] r_W_DATA; // @[AxiWrite.scala 83:33:@43692.4]
  reg [31:0] _RAND_14;
  reg  r_W_LAST; // @[AxiWrite.scala 84:33:@43693.4]
  reg [31:0] _RAND_15;
  reg [3:0] r_W_STRB; // @[AxiWrite.scala 85:33:@43694.4]
  reg [31:0] _RAND_16;
  reg  r_W_VALID; // @[AxiWrite.scala 86:33:@43695.4]
  reg [31:0] _RAND_17;
  reg  r_W_ID; // @[AxiWrite.scala 87:33:@43696.4]
  reg [31:0] _RAND_18;
  reg  r_B_READY; // @[AxiWrite.scala 90:33:@43697.4]
  reg [31:0] _RAND_19;
  reg [2:0] r_transaction_cnt; // @[AxiWrite.scala 93:44:@43698.4]
  reg [31:0] _RAND_20;
  reg [7:0] r_len; // @[AxiWrite.scala 94:44:@43699.4]
  reg [31:0] _RAND_21;
  wire [1:0] _T_192; // @[AxiWrite.scala 99:45:@43702.4]
  wire [1:0] _GEN_116; // @[AxiWrite.scala 99:43:@43703.4]
  wire [1:0] _T_193; // @[AxiWrite.scala 99:43:@43703.4]
  reg [1:0] state; // @[AxiWrite.scala 108:28:@43705.4]
  reg [31:0] _RAND_22;
  wire  _T_195; // @[Conditional.scala 37:30:@43706.4]
  wire  _T_199; // @[AxiWrite.scala 115:45:@43710.8]
  wire [3:0] _T_219; // @[AxiWrite.scala 145:68:@43736.12]
  wire [2:0] _T_220; // @[AxiWrite.scala 145:68:@43737.12]
  wire [2:0] _GEN_2; // @[AxiWrite.scala 140:50:@43730.10]
  wire [1:0] _GEN_3; // @[AxiWrite.scala 140:50:@43730.10]
  wire  _GEN_4; // @[AxiWrite.scala 140:50:@43730.10]
  wire  _GEN_13; // @[AxiWrite.scala 148:50:@43743.10]
  wire [2:0] _GEN_14; // @[AxiWrite.scala 148:50:@43743.10]
  wire  _GEN_15; // @[AxiWrite.scala 115:53:@43711.8]
  wire [7:0] _GEN_16; // @[AxiWrite.scala 115:53:@43711.8]
  wire [2:0] _GEN_17; // @[AxiWrite.scala 115:53:@43711.8]
  wire [1:0] _GEN_18; // @[AxiWrite.scala 115:53:@43711.8]
  wire  _GEN_19; // @[AxiWrite.scala 115:53:@43711.8]
  wire [3:0] _GEN_20; // @[AxiWrite.scala 115:53:@43711.8]
  wire [2:0] _GEN_21; // @[AxiWrite.scala 115:53:@43711.8]
  wire [3:0] _GEN_22; // @[AxiWrite.scala 115:53:@43711.8]
  wire [3:0] _GEN_23; // @[AxiWrite.scala 115:53:@43711.8]
  wire  _GEN_24; // @[AxiWrite.scala 115:53:@43711.8]
  wire [30:0] _GEN_25; // @[AxiWrite.scala 115:53:@43711.8]
  wire [7:0] _GEN_26; // @[AxiWrite.scala 115:53:@43711.8]
  wire  _GEN_27; // @[AxiWrite.scala 115:53:@43711.8]
  wire [31:0] _GEN_28; // @[AxiWrite.scala 115:53:@43711.8]
  wire [3:0] _GEN_29; // @[AxiWrite.scala 115:53:@43711.8]
  wire  _GEN_30; // @[AxiWrite.scala 115:53:@43711.8]
  wire [2:0] _GEN_32; // @[AxiWrite.scala 115:53:@43711.8]
  wire [1:0] _GEN_33; // @[AxiWrite.scala 115:53:@43711.8]
  wire  _GEN_34; // @[AxiWrite.scala 114:56:@43709.6]
  wire [7:0] _GEN_35; // @[AxiWrite.scala 114:56:@43709.6]
  wire [2:0] _GEN_36; // @[AxiWrite.scala 114:56:@43709.6]
  wire [1:0] _GEN_37; // @[AxiWrite.scala 114:56:@43709.6]
  wire  _GEN_38; // @[AxiWrite.scala 114:56:@43709.6]
  wire [3:0] _GEN_39; // @[AxiWrite.scala 114:56:@43709.6]
  wire [2:0] _GEN_40; // @[AxiWrite.scala 114:56:@43709.6]
  wire [3:0] _GEN_41; // @[AxiWrite.scala 114:56:@43709.6]
  wire [3:0] _GEN_42; // @[AxiWrite.scala 114:56:@43709.6]
  wire  _GEN_43; // @[AxiWrite.scala 114:56:@43709.6]
  wire [30:0] _GEN_44; // @[AxiWrite.scala 114:56:@43709.6]
  wire [7:0] _GEN_45; // @[AxiWrite.scala 114:56:@43709.6]
  wire  _GEN_46; // @[AxiWrite.scala 114:56:@43709.6]
  wire [31:0] _GEN_47; // @[AxiWrite.scala 114:56:@43709.6]
  wire [3:0] _GEN_48; // @[AxiWrite.scala 114:56:@43709.6]
  wire  _GEN_49; // @[AxiWrite.scala 114:56:@43709.6]
  wire  _GEN_50; // @[AxiWrite.scala 114:56:@43709.6]
  wire [2:0] _GEN_51; // @[AxiWrite.scala 114:56:@43709.6]
  wire [1:0] _GEN_52; // @[AxiWrite.scala 114:56:@43709.6]
  wire  _T_231; // @[Conditional.scala 37:30:@43768.6]
  wire  _T_235; // @[AxiWrite.scala 171:33:@43772.10]
  wire [8:0] _T_237; // @[AxiWrite.scala 172:45:@43774.12]
  wire [8:0] _T_238; // @[AxiWrite.scala 172:45:@43775.12]
  wire [7:0] _T_239; // @[AxiWrite.scala 172:45:@43776.12]
  wire  _T_244; // @[AxiWrite.scala 177:37:@43784.12]
  wire  _GEN_53; // @[AxiWrite.scala 177:45:@43785.12]
  wire [7:0] _GEN_54; // @[AxiWrite.scala 171:40:@43773.10]
  wire [31:0] _GEN_55; // @[AxiWrite.scala 171:40:@43773.10]
  wire  _GEN_56; // @[AxiWrite.scala 171:40:@43773.10]
  wire [1:0] _GEN_57; // @[AxiWrite.scala 171:40:@43773.10]
  wire [2:0] _GEN_58; // @[AxiWrite.scala 171:40:@43773.10]
  wire  _GEN_59; // @[AxiWrite.scala 171:40:@43773.10]
  wire [3:0] _GEN_60; // @[AxiWrite.scala 171:40:@43773.10]
  wire  _GEN_61; // @[AxiWrite.scala 171:40:@43773.10]
  wire [7:0] _GEN_63; // @[AxiWrite.scala 170:41:@43771.8]
  wire [31:0] _GEN_64; // @[AxiWrite.scala 170:41:@43771.8]
  wire  _GEN_65; // @[AxiWrite.scala 170:41:@43771.8]
  wire [1:0] _GEN_66; // @[AxiWrite.scala 170:41:@43771.8]
  wire [2:0] _GEN_67; // @[AxiWrite.scala 170:41:@43771.8]
  wire  _GEN_68; // @[AxiWrite.scala 170:41:@43771.8]
  wire [3:0] _GEN_69; // @[AxiWrite.scala 170:41:@43771.8]
  wire  _GEN_70; // @[AxiWrite.scala 170:41:@43771.8]
  wire  _T_253; // @[Conditional.scala 37:30:@43813.8]
  wire  write_response_ready; // @[AxiWrite.scala 95:41:@43700.4 AxiWrite.scala 98:30:@43701.4 AxiWrite.scala 99:30:@43704.4]
  wire [1:0] _GEN_71; // @[AxiWrite.scala 202:53:@43817.10]
  wire  _GEN_72; // @[Conditional.scala 39:67:@43814.8]
  wire [1:0] _GEN_73; // @[Conditional.scala 39:67:@43814.8]
  wire [7:0] _GEN_74; // @[Conditional.scala 39:67:@43769.6]
  wire [31:0] _GEN_75; // @[Conditional.scala 39:67:@43769.6]
  wire  _GEN_76; // @[Conditional.scala 39:67:@43769.6]
  wire [1:0] _GEN_77; // @[Conditional.scala 39:67:@43769.6]
  wire [2:0] _GEN_78; // @[Conditional.scala 39:67:@43769.6]
  wire  _GEN_79; // @[Conditional.scala 39:67:@43769.6]
  wire [3:0] _GEN_80; // @[Conditional.scala 39:67:@43769.6]
  wire  _GEN_81; // @[Conditional.scala 39:67:@43769.6]
  wire  _GEN_82; // @[Conditional.scala 39:67:@43769.6]
  wire  _GEN_83; // @[Conditional.scala 40:58:@43707.4]
  wire [7:0] _GEN_84; // @[Conditional.scala 40:58:@43707.4]
  wire [2:0] _GEN_85; // @[Conditional.scala 40:58:@43707.4]
  wire [1:0] _GEN_86; // @[Conditional.scala 40:58:@43707.4]
  wire  _GEN_87; // @[Conditional.scala 40:58:@43707.4]
  wire [3:0] _GEN_88; // @[Conditional.scala 40:58:@43707.4]
  wire [2:0] _GEN_89; // @[Conditional.scala 40:58:@43707.4]
  wire [3:0] _GEN_90; // @[Conditional.scala 40:58:@43707.4]
  wire [3:0] _GEN_91; // @[Conditional.scala 40:58:@43707.4]
  wire  _GEN_92; // @[Conditional.scala 40:58:@43707.4]
  wire [30:0] _GEN_93; // @[Conditional.scala 40:58:@43707.4]
  wire [7:0] _GEN_94; // @[Conditional.scala 40:58:@43707.4]
  wire  _GEN_95; // @[Conditional.scala 40:58:@43707.4]
  wire [31:0] _GEN_96; // @[Conditional.scala 40:58:@43707.4]
  wire [3:0] _GEN_97; // @[Conditional.scala 40:58:@43707.4]
  wire  _GEN_98; // @[Conditional.scala 40:58:@43707.4]
  wire [2:0] _GEN_100; // @[Conditional.scala 40:58:@43707.4]
  wire [1:0] _GEN_101; // @[Conditional.scala 40:58:@43707.4]
  wire  _GEN_102; // @[Conditional.scala 40:58:@43707.4]
  wire  _GEN_103; // @[Conditional.scala 40:58:@43707.4]
  wire  _T_258; // @[AxiWrite.scala 210:20:@43821.4]
  wire  _T_259; // @[AxiWrite.scala 210:37:@43822.4]
  wire [3:0] _GEN_104; // @[AxiWrite.scala 212:36:@43825.6]
  wire [3:0] _GEN_105; // @[AxiWrite.scala 212:36:@43825.6]
  wire  _T_265; // @[AxiWrite.scala 213:26:@43828.6]
  wire  _GEN_106; // @[AxiWrite.scala 213:38:@43829.6]
  wire  _GEN_107; // @[AxiWrite.scala 210:66:@43823.4]
  wire [3:0] _GEN_108; // @[AxiWrite.scala 210:66:@43823.4]
  wire [3:0] _GEN_109; // @[AxiWrite.scala 210:66:@43823.4]
  wire  _T_269; // @[AxiWrite.scala 210:37:@43833.4]
  wire [3:0] _GEN_110; // @[AxiWrite.scala 212:36:@43836.6]
  wire [3:0] _GEN_111; // @[AxiWrite.scala 212:36:@43836.6]
  wire [3:0] _GEN_114; // @[AxiWrite.scala 210:66:@43834.4]
  wire [3:0] _GEN_115; // @[AxiWrite.scala 210:66:@43834.4]
  assign _T_126 = waitingForResponse_0 == 1'h0; // @[AxiWrite.scala 59:81:@43666.4]
  assign firstFreeIdx = _T_126 ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@43671.4]
  assign _T_146 = io_BRESP == 2'h0; // @[AxiWrite.scala 63:62:@43676.4]
  assign _T_192 = ~ io_BRESP; // @[AxiWrite.scala 99:45:@43702.4]
  assign _GEN_116 = {{1'd0}, io_BVALID}; // @[AxiWrite.scala 99:43:@43703.4]
  assign _T_193 = _GEN_116 & _T_192; // @[AxiWrite.scala 99:43:@43703.4]
  assign _T_195 = 2'h0 == state; // @[Conditional.scala 37:30:@43706.4]
  assign _T_199 = r_transaction_cnt == 3'h0; // @[AxiWrite.scala 115:45:@43710.8]
  assign _T_219 = r_transaction_cnt + 3'h1; // @[AxiWrite.scala 145:68:@43736.12]
  assign _T_220 = r_transaction_cnt + 3'h1; // @[AxiWrite.scala 145:68:@43737.12]
  assign _GEN_2 = io_AWREADY ? 3'h0 : _T_220; // @[AxiWrite.scala 140:50:@43730.10]
  assign _GEN_3 = io_AWREADY ? 2'h1 : state; // @[AxiWrite.scala 140:50:@43730.10]
  assign _GEN_4 = io_AWREADY ? 1'h0 : 1'h1; // @[AxiWrite.scala 140:50:@43730.10]
  assign _GEN_13 = io_AWREADY ? r_AW_ID : 1'h0; // @[AxiWrite.scala 148:50:@43743.10]
  assign _GEN_14 = io_AWREADY ? r_AW_PROT : 3'h0; // @[AxiWrite.scala 148:50:@43743.10]
  assign _GEN_15 = _T_199 ? 1'h0 : r_B_READY; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_16 = _T_199 ? 8'h0 : r_AW_LEN; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_17 = _T_199 ? 3'h5 : r_AW_SIZE; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_18 = _T_199 ? 2'h1 : r_AW_BURST; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_19 = _T_199 ? 1'h0 : r_AW_LOCK; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_20 = _T_199 ? 4'h0 : r_AW_CACHE; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_21 = _T_199 ? 3'h0 : _GEN_14; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_22 = _T_199 ? 4'h0 : r_AW_QOS; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_23 = _T_199 ? 4'h0 : r_AW_REGION; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_24 = _T_199 ? firstFreeIdx : _GEN_13; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_25 = _T_199 ? io_storeAddrToMem : {{25'd0}, r_AW_ADDR}; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_26 = _T_199 ? 8'h1 : r_len; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_27 = _T_199 ? _GEN_4 : _GEN_4; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_28 = _T_199 ? io_storeDataToMem : r_W_DATA; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_29 = _T_199 ? 4'hf : r_W_STRB; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_30 = _T_199 ? 1'h1 : r_W_VALID; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_32 = _T_199 ? _GEN_2 : _GEN_2; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_33 = _T_199 ? _GEN_3 : _GEN_3; // @[AxiWrite.scala 115:53:@43711.8]
  assign _GEN_34 = io_storeQIdxInToAW_valid ? _GEN_15 : r_B_READY; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_35 = io_storeQIdxInToAW_valid ? _GEN_16 : r_AW_LEN; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_36 = io_storeQIdxInToAW_valid ? _GEN_17 : r_AW_SIZE; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_37 = io_storeQIdxInToAW_valid ? _GEN_18 : r_AW_BURST; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_38 = io_storeQIdxInToAW_valid ? _GEN_19 : r_AW_LOCK; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_39 = io_storeQIdxInToAW_valid ? _GEN_20 : r_AW_CACHE; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_40 = io_storeQIdxInToAW_valid ? _GEN_21 : r_AW_PROT; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_41 = io_storeQIdxInToAW_valid ? _GEN_22 : r_AW_QOS; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_42 = io_storeQIdxInToAW_valid ? _GEN_23 : r_AW_REGION; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_43 = io_storeQIdxInToAW_valid ? _GEN_24 : r_AW_ID; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_44 = io_storeQIdxInToAW_valid ? _GEN_25 : {{25'd0}, r_AW_ADDR}; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_45 = io_storeQIdxInToAW_valid ? _GEN_26 : r_len; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_46 = io_storeQIdxInToAW_valid ? _GEN_27 : r_AW_VALID; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_47 = io_storeQIdxInToAW_valid ? _GEN_28 : r_W_DATA; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_48 = io_storeQIdxInToAW_valid ? _GEN_29 : r_W_STRB; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_49 = io_storeQIdxInToAW_valid ? _GEN_30 : r_W_VALID; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_50 = io_storeQIdxInToAW_valid ? _T_199 : 1'h0; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_51 = io_storeQIdxInToAW_valid ? _GEN_32 : r_transaction_cnt; // @[AxiWrite.scala 114:56:@43709.6]
  assign _GEN_52 = io_storeQIdxInToAW_valid ? _GEN_33 : 2'h0; // @[AxiWrite.scala 114:56:@43709.6]
  assign _T_231 = 2'h1 == state; // @[Conditional.scala 37:30:@43768.6]
  assign _T_235 = r_len > 8'h0; // @[AxiWrite.scala 171:33:@43772.10]
  assign _T_237 = r_len - 8'h1; // @[AxiWrite.scala 172:45:@43774.12]
  assign _T_238 = $unsigned(_T_237); // @[AxiWrite.scala 172:45:@43775.12]
  assign _T_239 = _T_238[7:0]; // @[AxiWrite.scala 172:45:@43776.12]
  assign _T_244 = r_len == 8'h1; // @[AxiWrite.scala 177:37:@43784.12]
  assign _GEN_53 = _T_244 ? 1'h1 : r_W_LAST; // @[AxiWrite.scala 177:45:@43785.12]
  assign _GEN_54 = _T_235 ? _T_239 : r_len; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_55 = _T_235 ? io_storeDataToMem : 32'h0; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_56 = _T_235 ? firstFreeIdx : r_W_ID; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_57 = _T_235 ? 2'h1 : 2'h2; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_58 = _T_235 ? _T_220 : 3'h0; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_59 = _T_235 ? _GEN_53 : 1'h0; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_60 = _T_235 ? r_W_STRB : 4'h0; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_61 = _T_235 ? r_W_VALID : 1'h0; // @[AxiWrite.scala 171:40:@43773.10]
  assign _GEN_63 = io_WREADY ? _GEN_54 : r_len; // @[AxiWrite.scala 170:41:@43771.8]
  assign _GEN_64 = io_WREADY ? _GEN_55 : _GEN_28; // @[AxiWrite.scala 170:41:@43771.8]
  assign _GEN_65 = io_WREADY ? _GEN_56 : r_W_ID; // @[AxiWrite.scala 170:41:@43771.8]
  assign _GEN_66 = io_WREADY ? _GEN_57 : 2'h1; // @[AxiWrite.scala 170:41:@43771.8]
  assign _GEN_67 = io_WREADY ? _GEN_58 : r_transaction_cnt; // @[AxiWrite.scala 170:41:@43771.8]
  assign _GEN_68 = io_WREADY ? _GEN_59 : r_W_LAST; // @[AxiWrite.scala 170:41:@43771.8]
  assign _GEN_69 = io_WREADY ? _GEN_60 : r_W_STRB; // @[AxiWrite.scala 170:41:@43771.8]
  assign _GEN_70 = io_WREADY ? _GEN_61 : r_W_VALID; // @[AxiWrite.scala 170:41:@43771.8]
  assign _T_253 = 2'h2 == state; // @[Conditional.scala 37:30:@43813.8]
  assign write_response_ready = _T_193[0]; // @[AxiWrite.scala 95:41:@43700.4 AxiWrite.scala 98:30:@43701.4 AxiWrite.scala 99:30:@43704.4]
  assign _GEN_71 = write_response_ready ? 2'h0 : state; // @[AxiWrite.scala 202:53:@43817.10]
  assign _GEN_72 = _T_253 ? 1'h1 : r_B_READY; // @[Conditional.scala 39:67:@43814.8]
  assign _GEN_73 = _T_253 ? _GEN_71 : state; // @[Conditional.scala 39:67:@43814.8]
  assign _GEN_74 = _T_231 ? _GEN_63 : r_len; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_75 = _T_231 ? _GEN_64 : r_W_DATA; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_76 = _T_231 ? _GEN_65 : r_W_ID; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_77 = _T_231 ? _GEN_66 : _GEN_73; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_78 = _T_231 ? _GEN_67 : r_transaction_cnt; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_79 = _T_231 ? _GEN_68 : r_W_LAST; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_80 = _T_231 ? _GEN_69 : r_W_STRB; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_81 = _T_231 ? _GEN_70 : r_W_VALID; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_82 = _T_231 ? r_B_READY : _GEN_72; // @[Conditional.scala 39:67:@43769.6]
  assign _GEN_83 = _T_195 ? _GEN_34 : _GEN_82; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_84 = _T_195 ? _GEN_35 : r_AW_LEN; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_85 = _T_195 ? _GEN_36 : r_AW_SIZE; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_86 = _T_195 ? _GEN_37 : r_AW_BURST; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_87 = _T_195 ? _GEN_38 : r_AW_LOCK; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_88 = _T_195 ? _GEN_39 : r_AW_CACHE; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_89 = _T_195 ? _GEN_40 : r_AW_PROT; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_90 = _T_195 ? _GEN_41 : r_AW_QOS; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_91 = _T_195 ? _GEN_42 : r_AW_REGION; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_92 = _T_195 ? _GEN_43 : r_AW_ID; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_93 = _T_195 ? _GEN_44 : {{25'd0}, r_AW_ADDR}; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_94 = _T_195 ? _GEN_45 : _GEN_74; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_95 = _T_195 ? _GEN_46 : r_AW_VALID; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_96 = _T_195 ? _GEN_47 : _GEN_75; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_97 = _T_195 ? _GEN_48 : _GEN_80; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_98 = _T_195 ? _GEN_49 : _GEN_81; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_100 = _T_195 ? _GEN_51 : _GEN_78; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_101 = _T_195 ? _GEN_52 : _GEN_77; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_102 = _T_195 ? r_W_ID : _GEN_76; // @[Conditional.scala 40:58:@43707.4]
  assign _GEN_103 = _T_195 ? r_W_LAST : _GEN_79; // @[Conditional.scala 40:58:@43707.4]
  assign _T_258 = 1'h0 == firstFreeIdx; // @[AxiWrite.scala 210:20:@43821.4]
  assign _T_259 = _T_258 & io_storeQIdxInToAW_ready; // @[AxiWrite.scala 210:37:@43822.4]
  assign _GEN_104 = 1'h0 == firstFreeIdx ? io_storeQIdxInToAW_bits : idxArray_0; // @[AxiWrite.scala 212:36:@43825.6]
  assign _GEN_105 = firstFreeIdx ? io_storeQIdxInToAW_bits : idxArray_1; // @[AxiWrite.scala 212:36:@43825.6]
  assign _T_265 = 1'h0 == io_BID; // @[AxiWrite.scala 213:26:@43828.6]
  assign _GEN_106 = _T_265 ? 1'h0 : waitingForResponse_0; // @[AxiWrite.scala 213:38:@43829.6]
  assign _GEN_107 = _T_259 ? 1'h1 : _GEN_106; // @[AxiWrite.scala 210:66:@43823.4]
  assign _GEN_108 = _T_259 ? _GEN_104 : idxArray_0; // @[AxiWrite.scala 210:66:@43823.4]
  assign _GEN_109 = _T_259 ? _GEN_105 : idxArray_1; // @[AxiWrite.scala 210:66:@43823.4]
  assign _T_269 = firstFreeIdx & io_storeQIdxInToAW_ready; // @[AxiWrite.scala 210:37:@43833.4]
  assign _GEN_110 = 1'h0 == firstFreeIdx ? io_storeQIdxInToAW_bits : _GEN_108; // @[AxiWrite.scala 212:36:@43836.6]
  assign _GEN_111 = firstFreeIdx ? io_storeQIdxInToAW_bits : _GEN_109; // @[AxiWrite.scala 212:36:@43836.6]
  assign _GEN_114 = _T_269 ? _GEN_110 : _GEN_108; // @[AxiWrite.scala 210:66:@43834.4]
  assign _GEN_115 = _T_269 ? _GEN_111 : _GEN_109; // @[AxiWrite.scala 210:66:@43834.4]
  assign io_storeQIdxInToAW_ready = _T_195 ? _GEN_50 : 1'h0; // @[AxiWrite.scala 65:34:@43680.4 AxiWrite.scala 138:50:@43728.10]
  assign io_storeQIdxOutFromAW = io_BID ? idxArray_1 : idxArray_0; // @[AxiWrite.scala 64:36:@43679.4]
  assign io_storeQIdxOutFromAWValid = io_BVALID & _T_146; // @[AxiWrite.scala 63:36:@43678.4]
  assign io_AWID = r_AW_ID; // @[AxiWrite.scala 225:20:@43847.4]
  assign io_AWADDR = {{25'd0}, r_AW_ADDR}; // @[AxiWrite.scala 222:20:@43844.4]
  assign io_AWLEN = r_AW_LEN; // @[AxiWrite.scala 223:20:@43845.4]
  assign io_AWSIZE = r_AW_SIZE; // @[AxiWrite.scala 224:20:@43846.4]
  assign io_AWBURST = r_AW_BURST; // @[AxiWrite.scala 221:20:@43843.4]
  assign io_AWPROT = r_AW_PROT; // @[AxiWrite.scala 227:20:@43850.4]
  assign io_AWVALID = r_AW_VALID; // @[AxiWrite.scala 226:20:@43849.4]
  assign io_AWLOCK = r_AW_LOCK; // @[AxiWrite.scala 230:20:@43854.4]
  assign io_AWCACHE = r_AW_CACHE; // @[AxiWrite.scala 231:20:@43855.4]
  assign io_AWQOS = r_AW_QOS; // @[AxiWrite.scala 228:20:@43851.4]
  assign io_AWREGION = r_AW_REGION; // @[AxiWrite.scala 229:21:@43852.4]
  assign io_WID = r_W_ID; // @[AxiWrite.scala 238:20:@43862.4]
  assign io_WDATA = r_W_DATA; // @[AxiWrite.scala 234:20:@43856.4]
  assign io_WSTRB = r_W_STRB; // @[AxiWrite.scala 236:20:@43859.4]
  assign io_WLAST = r_W_LAST; // @[AxiWrite.scala 235:20:@43858.4]
  assign io_WVALID = r_W_VALID; // @[AxiWrite.scala 237:20:@43861.4]
  assign io_BREADY = r_B_READY; // @[AxiWrite.scala 241:20:@43864.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  idxArray_0 = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  idxArray_1 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  waitingForResponse_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  r_AW_BURST = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  r_AW_ADDR = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  r_AW_LEN = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  r_AW_SIZE = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  r_AW_ID = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  r_AW_VALID = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  r_AW_PROT = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  r_AW_QOS = _RAND_10[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  r_AW_LOCK = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  r_AW_CACHE = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  r_AW_REGION = _RAND_13[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  r_W_DATA = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  r_W_LAST = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_W_STRB = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  r_W_VALID = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  r_W_ID = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  r_B_READY = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  r_transaction_cnt = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  r_len = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  state = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      idxArray_0 <= 4'h0;
    end else begin
      if (_T_269) begin
        if (1'h0 == firstFreeIdx) begin
          idxArray_0 <= io_storeQIdxInToAW_bits;
        end else begin
          if (_T_259) begin
            if (1'h0 == firstFreeIdx) begin
              idxArray_0 <= io_storeQIdxInToAW_bits;
            end
          end
        end
      end else begin
        if (_T_259) begin
          if (1'h0 == firstFreeIdx) begin
            idxArray_0 <= io_storeQIdxInToAW_bits;
          end
        end
      end
    end
    if (reset) begin
      idxArray_1 <= 4'h0;
    end else begin
      if (_T_269) begin
        if (firstFreeIdx) begin
          idxArray_1 <= io_storeQIdxInToAW_bits;
        end else begin
          if (_T_259) begin
            if (firstFreeIdx) begin
              idxArray_1 <= io_storeQIdxInToAW_bits;
            end
          end
        end
      end else begin
        if (_T_259) begin
          if (firstFreeIdx) begin
            idxArray_1 <= io_storeQIdxInToAW_bits;
          end
        end
      end
    end
    if (reset) begin
      waitingForResponse_0 <= 1'h0;
    end else begin
      if (_T_259) begin
        waitingForResponse_0 <= 1'h1;
      end else begin
        if (_T_265) begin
          waitingForResponse_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      r_AW_BURST <= 2'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_BURST <= 2'h1;
          end
        end
      end
    end
    if (reset) begin
      r_AW_ADDR <= 6'h0;
    end else begin
      r_AW_ADDR <= _GEN_93[5:0];
    end
    if (reset) begin
      r_AW_LEN <= 8'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_LEN <= 8'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AW_SIZE <= 3'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_SIZE <= 3'h5;
          end
        end
      end
    end
    if (reset) begin
      r_AW_ID <= 1'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            if (_T_126) begin
              r_AW_ID <= 1'h0;
            end else begin
              r_AW_ID <= 1'h1;
            end
          end else begin
            if (!(io_AWREADY)) begin
              r_AW_ID <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AW_VALID <= 1'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            if (io_AWREADY) begin
              r_AW_VALID <= 1'h0;
            end else begin
              r_AW_VALID <= 1'h1;
            end
          end else begin
            if (io_AWREADY) begin
              r_AW_VALID <= 1'h0;
            end else begin
              r_AW_VALID <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AW_PROT <= 3'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_PROT <= 3'h0;
          end else begin
            if (!(io_AWREADY)) begin
              r_AW_PROT <= 3'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AW_QOS <= 4'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_QOS <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AW_LOCK <= 1'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_LOCK <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AW_CACHE <= 4'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_CACHE <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AW_REGION <= 4'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_AW_REGION <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      r_W_DATA <= 32'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_W_DATA <= io_storeDataToMem;
          end
        end
      end else begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (_T_235) begin
              r_W_DATA <= io_storeDataToMem;
            end else begin
              r_W_DATA <= 32'h0;
            end
          end else begin
            if (_T_199) begin
              r_W_DATA <= io_storeDataToMem;
            end
          end
        end
      end
    end
    if (reset) begin
      r_W_LAST <= 1'h0;
    end else begin
      if (!(_T_195)) begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (_T_235) begin
              if (_T_244) begin
                r_W_LAST <= 1'h1;
              end
            end else begin
              r_W_LAST <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_W_STRB <= 4'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_W_STRB <= 4'hf;
          end
        end
      end else begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (!(_T_235)) begin
              r_W_STRB <= 4'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_W_VALID <= 1'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_W_VALID <= 1'h1;
          end
        end
      end else begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (!(_T_235)) begin
              r_W_VALID <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_W_ID <= 1'h0;
    end else begin
      if (!(_T_195)) begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (_T_235) begin
              if (_T_126) begin
                r_W_ID <= 1'h0;
              end else begin
                r_W_ID <= 1'h1;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      r_B_READY <= 1'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_B_READY <= 1'h0;
          end
        end
      end else begin
        if (!(_T_231)) begin
          if (_T_253) begin
            r_B_READY <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      r_transaction_cnt <= 3'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            if (io_AWREADY) begin
              r_transaction_cnt <= 3'h0;
            end else begin
              r_transaction_cnt <= _T_220;
            end
          end else begin
            if (io_AWREADY) begin
              r_transaction_cnt <= 3'h0;
            end else begin
              r_transaction_cnt <= _T_220;
            end
          end
        end
      end else begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (_T_235) begin
              r_transaction_cnt <= _T_220;
            end else begin
              r_transaction_cnt <= 3'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_len <= 8'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            r_len <= 8'h1;
          end
        end
      end else begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (_T_235) begin
              r_len <= _T_239;
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_195) begin
        if (io_storeQIdxInToAW_valid) begin
          if (_T_199) begin
            if (io_AWREADY) begin
              state <= 2'h1;
            end
          end else begin
            if (io_AWREADY) begin
              state <= 2'h1;
            end
          end
        end else begin
          state <= 2'h0;
        end
      end else begin
        if (_T_231) begin
          if (io_WREADY) begin
            if (_T_235) begin
              state <= 2'h1;
            end else begin
              state <= 2'h2;
            end
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_253) begin
            if (write_response_ready) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
  end
endmodule
module AXI_READ( // @[:@43866.2]
  input         clock, // @[:@43867.4]
  input         reset, // @[:@43868.4]
  output [31:0] io_loadDataFromMem, // @[:@43869.4]
  input  [30:0] io_loadAddrToMem, // @[:@43869.4]
  output [31:0] io_loadQIdxForDataOut, // @[:@43869.4]
  output        io_loadQIdxForDataOutValid, // @[:@43869.4]
  output        io_loadQIdxForAddrIn_ready, // @[:@43869.4]
  input         io_loadQIdxForAddrIn_valid, // @[:@43869.4]
  input  [30:0] io_loadQIdxForAddrIn_bits, // @[:@43869.4]
  output        io_ARID, // @[:@43869.4]
  output [30:0] io_ARADDR, // @[:@43869.4]
  output [7:0]  io_ARLEN, // @[:@43869.4]
  output [2:0]  io_ARSIZE, // @[:@43869.4]
  output [1:0]  io_ARBURST, // @[:@43869.4]
  output        io_ARLOCK, // @[:@43869.4]
  output [3:0]  io_ARCACHE, // @[:@43869.4]
  output [3:0]  io_ARQOS, // @[:@43869.4]
  output [3:0]  io_ARREGION, // @[:@43869.4]
  output [2:0]  io_ARPROT, // @[:@43869.4]
  output        io_ARVALID, // @[:@43869.4]
  input         io_ARREADY, // @[:@43869.4]
  input         io_RID, // @[:@43869.4]
  input  [31:0] io_RDATA, // @[:@43869.4]
  input  [1:0]  io_RRESP, // @[:@43869.4]
  input         io_RLAST, // @[:@43869.4]
  input         io_RVALID, // @[:@43869.4]
  output        io_RREADY // @[:@43869.4]
);
  reg  r_AR_ID; // @[AxiRead.scala 50:27:@43871.4]
  reg [31:0] _RAND_0;
  reg [30:0] r_AR_ADDR; // @[AxiRead.scala 51:27:@43872.4]
  reg [31:0] _RAND_1;
  reg [7:0] r_AR_LEN; // @[AxiRead.scala 52:27:@43873.4]
  reg [31:0] _RAND_2;
  reg [2:0] r_AR_SIZE; // @[AxiRead.scala 53:27:@43874.4]
  reg [31:0] _RAND_3;
  reg [1:0] r_AR_BURST; // @[AxiRead.scala 54:27:@43875.4]
  reg [31:0] _RAND_4;
  reg [3:0] r_AR_QOS; // @[AxiRead.scala 55:28:@43876.4]
  reg [31:0] _RAND_5;
  reg  r_AR_LOCK; // @[AxiRead.scala 56:28:@43877.4]
  reg [31:0] _RAND_6;
  reg [3:0] r_AR_CACHE; // @[AxiRead.scala 57:28:@43878.4]
  reg [31:0] _RAND_7;
  reg [3:0] r_AR_REGION; // @[AxiRead.scala 58:28:@43879.4]
  reg [31:0] _RAND_8;
  reg [2:0] r_AR_PROT; // @[AxiRead.scala 59:27:@43880.4]
  reg [31:0] _RAND_9;
  reg  r_AR_VALID; // @[AxiRead.scala 60:27:@43881.4]
  reg [31:0] _RAND_10;
  reg [31:0] r_R_RDATA; // @[AxiRead.scala 65:27:@43883.4]
  reg [31:0] _RAND_11;
  reg  r_R_READY; // @[AxiRead.scala 66:27:@43884.4]
  reg [31:0] _RAND_12;
  reg [2:0] rx_transaction_cnt; // @[AxiRead.scala 69:38:@43885.4]
  reg [31:0] _RAND_13;
  reg [7:0] rx_len; // @[AxiRead.scala 70:38:@43886.4]
  reg [31:0] _RAND_14;
  wire [1:0] _T_95; // @[AxiRead.scala 75:39:@43889.4]
  wire [1:0] _GEN_81; // @[AxiRead.scala 75:37:@43890.4]
  wire [1:0] _T_96; // @[AxiRead.scala 75:37:@43890.4]
  wire [1:0] _GEN_82; // @[AxiRead.scala 75:49:@43891.4]
  wire [1:0] _T_97; // @[AxiRead.scala 75:49:@43891.4]
  reg [3:0] idxArray_0; // @[AxiRead.scala 78:25:@43896.4]
  reg [31:0] _RAND_15;
  reg [3:0] idxArray_1; // @[AxiRead.scala 78:25:@43896.4]
  reg [31:0] _RAND_16;
  reg  waitingForData_0; // @[AxiRead.scala 79:31:@43900.4]
  reg [31:0] _RAND_17;
  reg  waitingForData_1; // @[AxiRead.scala 79:31:@43900.4]
  reg [31:0] _RAND_18;
  wire  _T_155; // @[AxiRead.scala 80:71:@43901.4]
  wire  _T_157; // @[AxiRead.scala 80:71:@43902.4]
  wire  firstFreeIdx; // @[Mux.scala 31:69:@43906.4]
  wire  hasFreeIdx; // @[AxiRead.scala 81:41:@43910.4]
  reg [1:0] rx_state; // @[AxiRead.scala 91:25:@43911.4]
  reg [31:0] _RAND_19;
  wire  _T_175; // @[Conditional.scala 37:30:@43912.4]
  wire  _T_179; // @[AxiRead.scala 97:41:@43916.8]
  wire  _T_189; // @[AxiRead.scala 109:46:@43928.10]
  wire [3:0] _T_196; // @[AxiRead.scala 119:66:@43939.12]
  wire [2:0] _T_197; // @[AxiRead.scala 119:66:@43940.12]
  wire [2:0] _GEN_0; // @[AxiRead.scala 114:46:@43933.10]
  wire [1:0] _GEN_1; // @[AxiRead.scala 114:46:@43933.10]
  wire  _GEN_2; // @[AxiRead.scala 114:46:@43933.10]
  wire  _GEN_4; // @[AxiRead.scala 123:45:@43946.10]
  wire [30:0] _GEN_6; // @[AxiRead.scala 123:45:@43946.10]
  wire [1:0] _GEN_7; // @[AxiRead.scala 123:45:@43946.10]
  wire [7:0] _GEN_8; // @[AxiRead.scala 123:45:@43946.10]
  wire [2:0] _GEN_9; // @[AxiRead.scala 123:45:@43946.10]
  wire  _GEN_10; // @[AxiRead.scala 123:45:@43946.10]
  wire  _GEN_11; // @[AxiRead.scala 123:45:@43946.10]
  wire [2:0] _GEN_12; // @[AxiRead.scala 123:45:@43946.10]
  wire [30:0] _GEN_13; // @[AxiRead.scala 97:50:@43917.8]
  wire [7:0] _GEN_14; // @[AxiRead.scala 97:50:@43917.8]
  wire [2:0] _GEN_15; // @[AxiRead.scala 97:50:@43917.8]
  wire [1:0] _GEN_16; // @[AxiRead.scala 97:50:@43917.8]
  wire [7:0] _GEN_17; // @[AxiRead.scala 97:50:@43917.8]
  wire  _GEN_18; // @[AxiRead.scala 97:50:@43917.8]
  wire [3:0] _GEN_19; // @[AxiRead.scala 97:50:@43917.8]
  wire [2:0] _GEN_20; // @[AxiRead.scala 97:50:@43917.8]
  wire [3:0] _GEN_21; // @[AxiRead.scala 97:50:@43917.8]
  wire [3:0] _GEN_22; // @[AxiRead.scala 97:50:@43917.8]
  wire  _GEN_23; // @[AxiRead.scala 97:50:@43917.8]
  wire  _GEN_24; // @[AxiRead.scala 97:50:@43917.8]
  wire  _GEN_25; // @[AxiRead.scala 97:50:@43917.8]
  wire [2:0] _GEN_26; // @[AxiRead.scala 97:50:@43917.8]
  wire [1:0] _GEN_27; // @[AxiRead.scala 97:50:@43917.8]
  wire [30:0] _GEN_28; // @[AxiRead.scala 96:54:@43915.6]
  wire [7:0] _GEN_29; // @[AxiRead.scala 96:54:@43915.6]
  wire [2:0] _GEN_30; // @[AxiRead.scala 96:54:@43915.6]
  wire [1:0] _GEN_31; // @[AxiRead.scala 96:54:@43915.6]
  wire [7:0] _GEN_32; // @[AxiRead.scala 96:54:@43915.6]
  wire  _GEN_33; // @[AxiRead.scala 96:54:@43915.6]
  wire [3:0] _GEN_34; // @[AxiRead.scala 96:54:@43915.6]
  wire [2:0] _GEN_35; // @[AxiRead.scala 96:54:@43915.6]
  wire [3:0] _GEN_36; // @[AxiRead.scala 96:54:@43915.6]
  wire [3:0] _GEN_37; // @[AxiRead.scala 96:54:@43915.6]
  wire  _GEN_38; // @[AxiRead.scala 96:54:@43915.6]
  wire  _GEN_39; // @[AxiRead.scala 96:54:@43915.6]
  wire  _GEN_40; // @[AxiRead.scala 96:54:@43915.6]
  wire [2:0] _GEN_41; // @[AxiRead.scala 96:54:@43915.6]
  wire [1:0] _GEN_42; // @[AxiRead.scala 96:54:@43915.6]
  wire  _T_212; // @[Conditional.scala 37:30:@43971.6]
  wire  _T_216; // @[AxiRead.scala 146:30:@43975.10]
  wire [8:0] _T_218; // @[AxiRead.scala 148:41:@43977.12]
  wire [8:0] _T_219; // @[AxiRead.scala 148:41:@43978.12]
  wire [7:0] _T_220; // @[AxiRead.scala 148:41:@43979.12]
  wire  read_response_ready; // @[AxiRead.scala 71:34:@43887.4 AxiRead.scala 74:24:@43888.4 AxiRead.scala 75:24:@43892.4]
  wire  _GEN_43; // @[AxiRead.scala 151:55:@43984.12]
  wire [1:0] _GEN_44; // @[AxiRead.scala 151:55:@43984.12]
  wire [7:0] _GEN_45; // @[AxiRead.scala 146:37:@43976.10]
  wire [31:0] _GEN_46; // @[AxiRead.scala 146:37:@43976.10]
  wire [1:0] _GEN_47; // @[AxiRead.scala 146:37:@43976.10]
  wire  _GEN_48; // @[AxiRead.scala 146:37:@43976.10]
  wire [7:0] _GEN_49; // @[AxiRead.scala 145:36:@43974.8]
  wire [31:0] _GEN_50; // @[AxiRead.scala 145:36:@43974.8]
  wire [1:0] _GEN_51; // @[AxiRead.scala 145:36:@43974.8]
  wire  _GEN_52; // @[AxiRead.scala 145:36:@43974.8]
  wire [7:0] _GEN_53; // @[Conditional.scala 39:67:@43972.6]
  wire [31:0] _GEN_54; // @[Conditional.scala 39:67:@43972.6]
  wire [1:0] _GEN_55; // @[Conditional.scala 39:67:@43972.6]
  wire  _GEN_56; // @[Conditional.scala 39:67:@43972.6]
  wire [30:0] _GEN_57; // @[Conditional.scala 40:58:@43913.4]
  wire [7:0] _GEN_58; // @[Conditional.scala 40:58:@43913.4]
  wire [2:0] _GEN_59; // @[Conditional.scala 40:58:@43913.4]
  wire [1:0] _GEN_60; // @[Conditional.scala 40:58:@43913.4]
  wire [7:0] _GEN_61; // @[Conditional.scala 40:58:@43913.4]
  wire  _GEN_62; // @[Conditional.scala 40:58:@43913.4]
  wire [3:0] _GEN_63; // @[Conditional.scala 40:58:@43913.4]
  wire [2:0] _GEN_64; // @[Conditional.scala 40:58:@43913.4]
  wire [3:0] _GEN_65; // @[Conditional.scala 40:58:@43913.4]
  wire [3:0] _GEN_66; // @[Conditional.scala 40:58:@43913.4]
  wire  _GEN_67; // @[Conditional.scala 40:58:@43913.4]
  wire  _GEN_68; // @[Conditional.scala 40:58:@43913.4]
  wire  _GEN_69; // @[Conditional.scala 40:58:@43913.4]
  wire [2:0] _GEN_70; // @[Conditional.scala 40:58:@43913.4]
  wire [1:0] _GEN_71; // @[Conditional.scala 40:58:@43913.4]
  wire [31:0] _GEN_72; // @[Conditional.scala 40:58:@43913.4]
  wire [3:0] _GEN_74; // @[AxiRead.scala 165:25:@43997.4]
  wire  _T_230; // @[AxiRead.scala 166:56:@43998.4]
  wire  _T_233; // @[AxiRead.scala 171:14:@44001.4]
  wire  _T_234; // @[AxiRead.scala 171:31:@44002.4]
  wire  _T_235; // @[AxiRead.scala 171:45:@44003.4]
  wire  _T_236; // @[AxiRead.scala 171:59:@44004.4]
  wire  _T_239; // @[AxiRead.scala 174:21:@44010.6]
  wire  _T_240; // @[AxiRead.scala 174:32:@44011.6]
  wire  _T_243; // @[AxiRead.scala 174:45:@44013.6]
  wire  _GEN_75; // @[AxiRead.scala 174:65:@44014.6]
  wire [30:0] _GEN_76; // @[AxiRead.scala 171:90:@44005.4]
  wire  _GEN_77; // @[AxiRead.scala 171:90:@44005.4]
  wire  _T_247; // @[AxiRead.scala 171:31:@44018.4]
  wire  _T_248; // @[AxiRead.scala 171:45:@44019.4]
  wire  _T_249; // @[AxiRead.scala 171:59:@44020.4]
  wire  _T_253; // @[AxiRead.scala 174:32:@44027.6]
  wire  _T_256; // @[AxiRead.scala 174:45:@44029.6]
  wire  _GEN_78; // @[AxiRead.scala 174:65:@44030.6]
  wire [30:0] _GEN_79; // @[AxiRead.scala 171:90:@44021.4]
  wire  _GEN_80; // @[AxiRead.scala 171:90:@44021.4]
  assign _T_95 = ~ io_RRESP; // @[AxiRead.scala 75:39:@43889.4]
  assign _GEN_81 = {{1'd0}, io_RVALID}; // @[AxiRead.scala 75:37:@43890.4]
  assign _T_96 = _GEN_81 & _T_95; // @[AxiRead.scala 75:37:@43890.4]
  assign _GEN_82 = {{1'd0}, io_RLAST}; // @[AxiRead.scala 75:49:@43891.4]
  assign _T_97 = _T_96 & _GEN_82; // @[AxiRead.scala 75:49:@43891.4]
  assign _T_155 = waitingForData_0 == 1'h0; // @[AxiRead.scala 80:71:@43901.4]
  assign _T_157 = waitingForData_1 == 1'h0; // @[AxiRead.scala 80:71:@43902.4]
  assign firstFreeIdx = _T_155 ? 1'h0 : 1'h1; // @[Mux.scala 31:69:@43906.4]
  assign hasFreeIdx = _T_155 | _T_157; // @[AxiRead.scala 81:41:@43910.4]
  assign _T_175 = 2'h0 == rx_state; // @[Conditional.scala 37:30:@43912.4]
  assign _T_179 = rx_transaction_cnt == 3'h0; // @[AxiRead.scala 97:41:@43916.8]
  assign _T_189 = hasFreeIdx & io_loadQIdxForAddrIn_valid; // @[AxiRead.scala 109:46:@43928.10]
  assign _T_196 = rx_transaction_cnt + 3'h1; // @[AxiRead.scala 119:66:@43939.12]
  assign _T_197 = rx_transaction_cnt + 3'h1; // @[AxiRead.scala 119:66:@43940.12]
  assign _GEN_0 = io_ARREADY ? 3'h0 : _T_197; // @[AxiRead.scala 114:46:@43933.10]
  assign _GEN_1 = io_ARREADY ? 2'h1 : rx_state; // @[AxiRead.scala 114:46:@43933.10]
  assign _GEN_2 = io_ARREADY ? 1'h0 : _T_189; // @[AxiRead.scala 114:46:@43933.10]
  assign _GEN_4 = io_ARREADY ? 1'h0 : 1'h1; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_6 = io_ARREADY ? r_AR_ADDR : io_loadAddrToMem; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_7 = io_ARREADY ? r_AR_BURST : 2'h1; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_8 = io_ARREADY ? r_AR_LEN : 8'h0; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_9 = io_ARREADY ? r_AR_SIZE : 3'h5; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_10 = io_ARREADY ? r_R_READY : 1'h1; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_11 = io_ARREADY ? r_AR_ID : 1'h0; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_12 = io_ARREADY ? r_AR_PROT : 3'h0; // @[AxiRead.scala 123:45:@43946.10]
  assign _GEN_13 = _T_179 ? io_loadAddrToMem : _GEN_6; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_14 = _T_179 ? 8'h0 : _GEN_8; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_15 = _T_179 ? 3'h5 : _GEN_9; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_16 = _T_179 ? 2'h1 : _GEN_7; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_17 = _T_179 ? 8'h1 : rx_len; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_18 = _T_179 ? 1'h0 : r_AR_LOCK; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_19 = _T_179 ? 4'h0 : r_AR_CACHE; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_20 = _T_179 ? 3'h0 : _GEN_12; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_21 = _T_179 ? 4'h0 : r_AR_QOS; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_22 = _T_179 ? 4'h0 : r_AR_REGION; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_23 = _T_179 ? _GEN_2 : _GEN_4; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_24 = _T_179 ? firstFreeIdx : _GEN_11; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_25 = _T_179 ? 1'h1 : _GEN_10; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_26 = _T_179 ? _GEN_0 : _GEN_0; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_27 = _T_179 ? _GEN_1 : _GEN_1; // @[AxiRead.scala 97:50:@43917.8]
  assign _GEN_28 = io_loadQIdxForAddrIn_valid ? _GEN_13 : r_AR_ADDR; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_29 = io_loadQIdxForAddrIn_valid ? _GEN_14 : r_AR_LEN; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_30 = io_loadQIdxForAddrIn_valid ? _GEN_15 : r_AR_SIZE; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_31 = io_loadQIdxForAddrIn_valid ? _GEN_16 : r_AR_BURST; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_32 = io_loadQIdxForAddrIn_valid ? _GEN_17 : rx_len; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_33 = io_loadQIdxForAddrIn_valid ? _GEN_18 : r_AR_LOCK; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_34 = io_loadQIdxForAddrIn_valid ? _GEN_19 : r_AR_CACHE; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_35 = io_loadQIdxForAddrIn_valid ? _GEN_20 : r_AR_PROT; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_36 = io_loadQIdxForAddrIn_valid ? _GEN_21 : r_AR_QOS; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_37 = io_loadQIdxForAddrIn_valid ? _GEN_22 : r_AR_REGION; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_38 = io_loadQIdxForAddrIn_valid ? _GEN_23 : r_AR_VALID; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_39 = io_loadQIdxForAddrIn_valid ? _GEN_24 : r_AR_ID; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_40 = io_loadQIdxForAddrIn_valid ? _GEN_25 : r_R_READY; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_41 = io_loadQIdxForAddrIn_valid ? _GEN_26 : rx_transaction_cnt; // @[AxiRead.scala 96:54:@43915.6]
  assign _GEN_42 = io_loadQIdxForAddrIn_valid ? _GEN_27 : 2'h0; // @[AxiRead.scala 96:54:@43915.6]
  assign _T_212 = 2'h1 == rx_state; // @[Conditional.scala 37:30:@43971.6]
  assign _T_216 = rx_len >= 8'h1; // @[AxiRead.scala 146:30:@43975.10]
  assign _T_218 = rx_len - 8'h1; // @[AxiRead.scala 148:41:@43977.12]
  assign _T_219 = $unsigned(_T_218); // @[AxiRead.scala 148:41:@43978.12]
  assign _T_220 = _T_219[7:0]; // @[AxiRead.scala 148:41:@43979.12]
  assign read_response_ready = _T_97[0]; // @[AxiRead.scala 71:34:@43887.4 AxiRead.scala 74:24:@43888.4 AxiRead.scala 75:24:@43892.4]
  assign _GEN_43 = read_response_ready ? 1'h0 : r_R_READY; // @[AxiRead.scala 151:55:@43984.12]
  assign _GEN_44 = read_response_ready ? 2'h0 : 2'h1; // @[AxiRead.scala 151:55:@43984.12]
  assign _GEN_45 = _T_216 ? _T_220 : rx_len; // @[AxiRead.scala 146:37:@43976.10]
  assign _GEN_46 = _T_216 ? io_RDATA : r_R_RDATA; // @[AxiRead.scala 146:37:@43976.10]
  assign _GEN_47 = _T_216 ? _GEN_44 : rx_state; // @[AxiRead.scala 146:37:@43976.10]
  assign _GEN_48 = _T_216 ? _GEN_43 : r_R_READY; // @[AxiRead.scala 146:37:@43976.10]
  assign _GEN_49 = io_RVALID ? _GEN_45 : rx_len; // @[AxiRead.scala 145:36:@43974.8]
  assign _GEN_50 = io_RVALID ? _GEN_46 : 32'h0; // @[AxiRead.scala 145:36:@43974.8]
  assign _GEN_51 = io_RVALID ? _GEN_47 : 2'h1; // @[AxiRead.scala 145:36:@43974.8]
  assign _GEN_52 = io_RVALID ? _GEN_48 : r_R_READY; // @[AxiRead.scala 145:36:@43974.8]
  assign _GEN_53 = _T_212 ? _GEN_49 : rx_len; // @[Conditional.scala 39:67:@43972.6]
  assign _GEN_54 = _T_212 ? _GEN_50 : r_R_RDATA; // @[Conditional.scala 39:67:@43972.6]
  assign _GEN_55 = _T_212 ? _GEN_51 : rx_state; // @[Conditional.scala 39:67:@43972.6]
  assign _GEN_56 = _T_212 ? _GEN_52 : r_R_READY; // @[Conditional.scala 39:67:@43972.6]
  assign _GEN_57 = _T_175 ? _GEN_28 : r_AR_ADDR; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_58 = _T_175 ? _GEN_29 : r_AR_LEN; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_59 = _T_175 ? _GEN_30 : r_AR_SIZE; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_60 = _T_175 ? _GEN_31 : r_AR_BURST; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_61 = _T_175 ? _GEN_32 : _GEN_53; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_62 = _T_175 ? _GEN_33 : r_AR_LOCK; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_63 = _T_175 ? _GEN_34 : r_AR_CACHE; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_64 = _T_175 ? _GEN_35 : r_AR_PROT; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_65 = _T_175 ? _GEN_36 : r_AR_QOS; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_66 = _T_175 ? _GEN_37 : r_AR_REGION; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_67 = _T_175 ? _GEN_38 : r_AR_VALID; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_68 = _T_175 ? _GEN_39 : r_AR_ID; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_69 = _T_175 ? _GEN_40 : _GEN_56; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_70 = _T_175 ? _GEN_41 : rx_transaction_cnt; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_71 = _T_175 ? _GEN_42 : _GEN_55; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_72 = _T_175 ? r_R_RDATA : _GEN_54; // @[Conditional.scala 40:58:@43913.4]
  assign _GEN_74 = io_RID ? idxArray_1 : idxArray_0; // @[AxiRead.scala 165:25:@43997.4]
  assign _T_230 = io_RRESP == 2'h0; // @[AxiRead.scala 166:56:@43998.4]
  assign _T_233 = 1'h0 == firstFreeIdx; // @[AxiRead.scala 171:14:@44001.4]
  assign _T_234 = _T_233 & hasFreeIdx; // @[AxiRead.scala 171:31:@44002.4]
  assign _T_235 = _T_234 & io_ARREADY; // @[AxiRead.scala 171:45:@44003.4]
  assign _T_236 = _T_235 & io_loadQIdxForAddrIn_valid; // @[AxiRead.scala 171:59:@44004.4]
  assign _T_239 = 1'h0 == io_RID; // @[AxiRead.scala 174:21:@44010.6]
  assign _T_240 = _T_239 & io_RVALID; // @[AxiRead.scala 174:32:@44011.6]
  assign _T_243 = _T_240 & _T_230; // @[AxiRead.scala 174:45:@44013.6]
  assign _GEN_75 = _T_243 ? 1'h0 : waitingForData_0; // @[AxiRead.scala 174:65:@44014.6]
  assign _GEN_76 = _T_236 ? io_loadQIdxForAddrIn_bits : {{27'd0}, idxArray_0}; // @[AxiRead.scala 171:90:@44005.4]
  assign _GEN_77 = _T_236 ? 1'h1 : _GEN_75; // @[AxiRead.scala 171:90:@44005.4]
  assign _T_247 = firstFreeIdx & hasFreeIdx; // @[AxiRead.scala 171:31:@44018.4]
  assign _T_248 = _T_247 & io_ARREADY; // @[AxiRead.scala 171:45:@44019.4]
  assign _T_249 = _T_248 & io_loadQIdxForAddrIn_valid; // @[AxiRead.scala 171:59:@44020.4]
  assign _T_253 = io_RID & io_RVALID; // @[AxiRead.scala 174:32:@44027.6]
  assign _T_256 = _T_253 & _T_230; // @[AxiRead.scala 174:45:@44029.6]
  assign _GEN_78 = _T_256 ? 1'h0 : waitingForData_1; // @[AxiRead.scala 174:65:@44030.6]
  assign _GEN_79 = _T_249 ? io_loadQIdxForAddrIn_bits : {{27'd0}, idxArray_1}; // @[AxiRead.scala 171:90:@44021.4]
  assign _GEN_80 = _T_249 ? 1'h1 : _GEN_78; // @[AxiRead.scala 171:90:@44021.4]
  assign io_loadDataFromMem = r_R_RDATA; // @[AxiRead.scala 198:24:@44048.4]
  assign io_loadQIdxForDataOut = {{28'd0}, _GEN_74}; // @[AxiRead.scala 165:25:@43997.4]
  assign io_loadQIdxForDataOutValid = io_RVALID & _T_230; // @[AxiRead.scala 166:30:@44000.4]
  assign io_loadQIdxForAddrIn_ready = hasFreeIdx & io_ARREADY; // @[AxiRead.scala 164:30:@43996.4]
  assign io_ARID = r_AR_ID; // @[AxiRead.scala 185:16:@44037.4]
  assign io_ARADDR = r_AR_ADDR; // @[AxiRead.scala 182:16:@44034.4]
  assign io_ARLEN = r_AR_LEN; // @[AxiRead.scala 183:16:@44035.4]
  assign io_ARSIZE = r_AR_SIZE; // @[AxiRead.scala 184:16:@44036.4]
  assign io_ARBURST = r_AR_BURST; // @[AxiRead.scala 181:16:@44033.4]
  assign io_ARLOCK = r_AR_LOCK; // @[AxiRead.scala 190:17:@44044.4]
  assign io_ARCACHE = r_AR_CACHE; // @[AxiRead.scala 191:17:@44045.4]
  assign io_ARQOS = r_AR_QOS; // @[AxiRead.scala 188:17:@44041.4]
  assign io_ARREGION = r_AR_REGION; // @[AxiRead.scala 189:17:@44042.4]
  assign io_ARPROT = r_AR_PROT; // @[AxiRead.scala 187:16:@44040.4]
  assign io_ARVALID = r_AR_VALID; // @[AxiRead.scala 186:16:@44039.4]
  assign io_RREADY = r_R_READY; // @[AxiRead.scala 194:17:@44047.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_AR_ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  r_AR_ADDR = _RAND_1[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  r_AR_LEN = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  r_AR_SIZE = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  r_AR_BURST = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  r_AR_QOS = _RAND_5[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  r_AR_LOCK = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  r_AR_CACHE = _RAND_7[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  r_AR_REGION = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  r_AR_PROT = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  r_AR_VALID = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  r_R_RDATA = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  r_R_READY = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  rx_transaction_cnt = _RAND_13[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  rx_len = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  idxArray_0 = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  idxArray_1 = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  waitingForData_0 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  waitingForData_1 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  rx_state = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      r_AR_ID <= 1'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            if (_T_155) begin
              r_AR_ID <= 1'h0;
            end else begin
              r_AR_ID <= 1'h1;
            end
          end else begin
            if (!(io_ARREADY)) begin
              r_AR_ID <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AR_ADDR <= 31'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_ADDR <= io_loadAddrToMem;
          end else begin
            if (!(io_ARREADY)) begin
              r_AR_ADDR <= io_loadAddrToMem;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AR_LEN <= 8'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_LEN <= 8'h0;
          end else begin
            if (!(io_ARREADY)) begin
              r_AR_LEN <= 8'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AR_SIZE <= 3'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_SIZE <= 3'h5;
          end else begin
            if (!(io_ARREADY)) begin
              r_AR_SIZE <= 3'h5;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AR_BURST <= 2'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_BURST <= 2'h1;
          end else begin
            if (!(io_ARREADY)) begin
              r_AR_BURST <= 2'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AR_QOS <= 4'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_QOS <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AR_LOCK <= 1'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_LOCK <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AR_CACHE <= 4'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_CACHE <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AR_REGION <= 4'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_REGION <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      r_AR_PROT <= 3'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_AR_PROT <= 3'h0;
          end else begin
            if (!(io_ARREADY)) begin
              r_AR_PROT <= 3'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      r_AR_VALID <= 1'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            if (io_ARREADY) begin
              r_AR_VALID <= 1'h0;
            end else begin
              r_AR_VALID <= _T_189;
            end
          end else begin
            if (io_ARREADY) begin
              r_AR_VALID <= 1'h0;
            end else begin
              r_AR_VALID <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      r_R_RDATA <= 32'h0;
    end else begin
      if (!(_T_175)) begin
        if (_T_212) begin
          if (io_RVALID) begin
            if (_T_216) begin
              r_R_RDATA <= io_RDATA;
            end
          end else begin
            r_R_RDATA <= 32'h0;
          end
        end
      end
    end
    if (reset) begin
      r_R_READY <= 1'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            r_R_READY <= 1'h1;
          end else begin
            if (!(io_ARREADY)) begin
              r_R_READY <= 1'h1;
            end
          end
        end
      end else begin
        if (_T_212) begin
          if (io_RVALID) begin
            if (_T_216) begin
              if (read_response_ready) begin
                r_R_READY <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      rx_transaction_cnt <= 3'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            if (io_ARREADY) begin
              rx_transaction_cnt <= 3'h0;
            end else begin
              rx_transaction_cnt <= _T_197;
            end
          end else begin
            if (io_ARREADY) begin
              rx_transaction_cnt <= 3'h0;
            end else begin
              rx_transaction_cnt <= _T_197;
            end
          end
        end
      end
    end
    if (reset) begin
      rx_len <= 8'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            rx_len <= 8'h1;
          end
        end
      end else begin
        if (_T_212) begin
          if (io_RVALID) begin
            if (_T_216) begin
              rx_len <= _T_220;
            end
          end
        end
      end
    end
    if (reset) begin
      idxArray_0 <= 4'h0;
    end else begin
      idxArray_0 <= _GEN_76[3:0];
    end
    if (reset) begin
      idxArray_1 <= 4'h0;
    end else begin
      idxArray_1 <= _GEN_79[3:0];
    end
    if (reset) begin
      waitingForData_0 <= 1'h0;
    end else begin
      if (_T_236) begin
        waitingForData_0 <= 1'h1;
      end else begin
        if (_T_243) begin
          waitingForData_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      waitingForData_1 <= 1'h0;
    end else begin
      if (_T_249) begin
        waitingForData_1 <= 1'h1;
      end else begin
        if (_T_256) begin
          waitingForData_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      rx_state <= 2'h0;
    end else begin
      if (_T_175) begin
        if (io_loadQIdxForAddrIn_valid) begin
          if (_T_179) begin
            if (io_ARREADY) begin
              rx_state <= 2'h1;
            end
          end else begin
            if (io_ARREADY) begin
              rx_state <= 2'h1;
            end
          end
        end else begin
          rx_state <= 2'h0;
        end
      end else begin
        if (_T_212) begin
          if (io_RVALID) begin
            if (_T_216) begin
              if (read_response_ready) begin
                rx_state <= 2'h0;
              end else begin
                rx_state <= 2'h1;
              end
            end
          end else begin
            rx_state <= 2'h1;
          end
        end
      end
    end
  end
endmodule
module LOAD_PORT_LSQ_a( // @[:@44050.2]
  input         clock, // @[:@44051.4]
  input         reset, // @[:@44052.4]
  output        io_addrFromPrev_ready, // @[:@44053.4]
  input         io_addrFromPrev_valid, // @[:@44053.4]
  input  [30:0] io_addrFromPrev_bits, // @[:@44053.4]
  input         io_portEnable, // @[:@44053.4]
  input         io_dataToNext_ready, // @[:@44053.4]
  output        io_dataToNext_valid, // @[:@44053.4]
  output [31:0] io_dataToNext_bits, // @[:@44053.4]
  output        io_loadAddrEnable, // @[:@44053.4]
  output [30:0] io_addrToLoadQueue, // @[:@44053.4]
  output        io_dataFromLoadQueue_ready, // @[:@44053.4]
  input         io_dataFromLoadQueue_valid, // @[:@44053.4]
  input  [31:0] io_dataFromLoadQueue_bits // @[:@44053.4]
);
  reg [4:0] cnt; // @[LoadPort.scala 23:20:@44055.4]
  reg [31:0] _RAND_0;
  wire  _T_44; // @[LoadPort.scala 26:25:@44056.4]
  wire  _T_45; // @[LoadPort.scala 26:22:@44057.4]
  wire  _T_47; // @[LoadPort.scala 26:51:@44058.4]
  wire  _T_48; // @[LoadPort.scala 26:44:@44059.4]
  wire [5:0] _T_50; // @[LoadPort.scala 27:16:@44061.6]
  wire [4:0] _T_51; // @[LoadPort.scala 27:16:@44062.6]
  wire  _T_53; // @[LoadPort.scala 28:35:@44066.6]
  wire  _T_54; // @[LoadPort.scala 28:32:@44067.6]
  wire  _T_56; // @[LoadPort.scala 28:57:@44068.6]
  wire  _T_57; // @[LoadPort.scala 28:50:@44069.6]
  wire [5:0] _T_59; // @[LoadPort.scala 29:16:@44071.8]
  wire [5:0] _T_60; // @[LoadPort.scala 29:16:@44072.8]
  wire [4:0] _T_61; // @[LoadPort.scala 29:16:@44073.8]
  wire [4:0] _GEN_0; // @[LoadPort.scala 28:66:@44070.6]
  wire [4:0] _GEN_1; // @[LoadPort.scala 26:75:@44060.4]
  wire  _T_63; // @[LoadPort.scala 33:28:@44077.4]
  assign _T_44 = io_loadAddrEnable == 1'h0; // @[LoadPort.scala 26:25:@44056.4]
  assign _T_45 = io_portEnable & _T_44; // @[LoadPort.scala 26:22:@44057.4]
  assign _T_47 = cnt != 5'h10; // @[LoadPort.scala 26:51:@44058.4]
  assign _T_48 = _T_45 & _T_47; // @[LoadPort.scala 26:44:@44059.4]
  assign _T_50 = cnt + 5'h1; // @[LoadPort.scala 27:16:@44061.6]
  assign _T_51 = cnt + 5'h1; // @[LoadPort.scala 27:16:@44062.6]
  assign _T_53 = io_portEnable == 1'h0; // @[LoadPort.scala 28:35:@44066.6]
  assign _T_54 = io_loadAddrEnable & _T_53; // @[LoadPort.scala 28:32:@44067.6]
  assign _T_56 = cnt != 5'h0; // @[LoadPort.scala 28:57:@44068.6]
  assign _T_57 = _T_54 & _T_56; // @[LoadPort.scala 28:50:@44069.6]
  assign _T_59 = cnt - 5'h1; // @[LoadPort.scala 29:16:@44071.8]
  assign _T_60 = $unsigned(_T_59); // @[LoadPort.scala 29:16:@44072.8]
  assign _T_61 = _T_60[4:0]; // @[LoadPort.scala 29:16:@44073.8]
  assign _GEN_0 = _T_57 ? _T_61 : cnt; // @[LoadPort.scala 28:66:@44070.6]
  assign _GEN_1 = _T_48 ? _T_51 : _GEN_0; // @[LoadPort.scala 26:75:@44060.4]
  assign _T_63 = cnt > 5'h0; // @[LoadPort.scala 33:28:@44077.4]
  assign io_addrFromPrev_ready = cnt > 5'h0; // @[LoadPort.scala 34:25:@44081.4]
  assign io_dataToNext_valid = io_dataFromLoadQueue_valid; // @[LoadPort.scala 35:17:@44083.4]
  assign io_dataToNext_bits = io_dataFromLoadQueue_bits; // @[LoadPort.scala 35:17:@44082.4]
  assign io_loadAddrEnable = _T_63 & io_addrFromPrev_valid; // @[LoadPort.scala 33:21:@44079.4]
  assign io_addrToLoadQueue = io_addrFromPrev_bits; // @[LoadPort.scala 32:22:@44076.4]
  assign io_dataFromLoadQueue_ready = io_dataToNext_ready; // @[LoadPort.scala 35:17:@44084.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_48) begin
        cnt <= _T_51;
      end else begin
        if (_T_57) begin
          cnt <= _T_61;
        end
      end
    end
  end
endmodule
module STORE_DATA_PORT_LSQ_a( // @[:@44086.2]
  input         clock, // @[:@44087.4]
  input         reset, // @[:@44088.4]
  output        io_dataFromPrev_ready, // @[:@44089.4]
  input         io_dataFromPrev_valid, // @[:@44089.4]
  input  [31:0] io_dataFromPrev_bits, // @[:@44089.4]
  input         io_portEnable, // @[:@44089.4]
  output        io_storeDataEnable, // @[:@44089.4]
  output [31:0] io_dataToStoreQueue // @[:@44089.4]
);
  reg [4:0] cnt; // @[StoreDataPort.scala 21:20:@44091.4]
  reg [31:0] _RAND_0;
  wire  _T_26; // @[StoreDataPort.scala 24:25:@44092.4]
  wire  _T_27; // @[StoreDataPort.scala 24:22:@44093.4]
  wire  _T_29; // @[StoreDataPort.scala 24:52:@44094.4]
  wire  _T_30; // @[StoreDataPort.scala 24:45:@44095.4]
  wire [5:0] _T_32; // @[StoreDataPort.scala 25:16:@44097.6]
  wire [4:0] _T_33; // @[StoreDataPort.scala 25:16:@44098.6]
  wire  _T_35; // @[StoreDataPort.scala 26:36:@44102.6]
  wire  _T_36; // @[StoreDataPort.scala 26:33:@44103.6]
  wire  _T_38; // @[StoreDataPort.scala 26:58:@44104.6]
  wire  _T_39; // @[StoreDataPort.scala 26:51:@44105.6]
  wire [5:0] _T_41; // @[StoreDataPort.scala 27:16:@44107.8]
  wire [5:0] _T_42; // @[StoreDataPort.scala 27:16:@44108.8]
  wire [4:0] _T_43; // @[StoreDataPort.scala 27:16:@44109.8]
  wire [4:0] _GEN_0; // @[StoreDataPort.scala 26:67:@44106.6]
  wire [4:0] _GEN_1; // @[StoreDataPort.scala 24:76:@44096.4]
  wire  _T_45; // @[StoreDataPort.scala 31:29:@44113.4]
  assign _T_26 = io_storeDataEnable == 1'h0; // @[StoreDataPort.scala 24:25:@44092.4]
  assign _T_27 = io_portEnable & _T_26; // @[StoreDataPort.scala 24:22:@44093.4]
  assign _T_29 = cnt != 5'h10; // @[StoreDataPort.scala 24:52:@44094.4]
  assign _T_30 = _T_27 & _T_29; // @[StoreDataPort.scala 24:45:@44095.4]
  assign _T_32 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@44097.6]
  assign _T_33 = cnt + 5'h1; // @[StoreDataPort.scala 25:16:@44098.6]
  assign _T_35 = io_portEnable == 1'h0; // @[StoreDataPort.scala 26:36:@44102.6]
  assign _T_36 = io_storeDataEnable & _T_35; // @[StoreDataPort.scala 26:33:@44103.6]
  assign _T_38 = cnt != 5'h0; // @[StoreDataPort.scala 26:58:@44104.6]
  assign _T_39 = _T_36 & _T_38; // @[StoreDataPort.scala 26:51:@44105.6]
  assign _T_41 = cnt - 5'h1; // @[StoreDataPort.scala 27:16:@44107.8]
  assign _T_42 = $unsigned(_T_41); // @[StoreDataPort.scala 27:16:@44108.8]
  assign _T_43 = _T_42[4:0]; // @[StoreDataPort.scala 27:16:@44109.8]
  assign _GEN_0 = _T_39 ? _T_43 : cnt; // @[StoreDataPort.scala 26:67:@44106.6]
  assign _GEN_1 = _T_30 ? _T_33 : _GEN_0; // @[StoreDataPort.scala 24:76:@44096.4]
  assign _T_45 = cnt > 5'h0; // @[StoreDataPort.scala 31:29:@44113.4]
  assign io_dataFromPrev_ready = cnt > 5'h0; // @[StoreDataPort.scala 32:25:@44117.4]
  assign io_storeDataEnable = _T_45 & io_dataFromPrev_valid; // @[StoreDataPort.scala 31:22:@44115.4]
  assign io_dataToStoreQueue = io_dataFromPrev_bits; // @[StoreDataPort.scala 30:23:@44112.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 5'h0;
    end else begin
      if (_T_30) begin
        cnt <= _T_33;
      end else begin
        if (_T_39) begin
          cnt <= _T_43;
        end
      end
    end
  end
endmodule
module LSQ_a( // @[:@44152.2]
  input         clock, // @[:@44153.4]
  input         reset, // @[:@44154.4]
  output        io_ARID, // @[:@44155.4]
  output [30:0] io_ARADDR, // @[:@44155.4]
  output [7:0]  io_ARLEN, // @[:@44155.4]
  output [2:0]  io_ARSIZE, // @[:@44155.4]
  output [1:0]  io_ARBURST, // @[:@44155.4]
  output        io_ARLOCK, // @[:@44155.4]
  output [3:0]  io_ARCACHE, // @[:@44155.4]
  output [2:0]  io_ARPROT, // @[:@44155.4]
  output [3:0]  io_ARQOS, // @[:@44155.4]
  output [3:0]  io_ARREGION, // @[:@44155.4]
  output        io_ARVALID, // @[:@44155.4]
  input         io_ARREADY, // @[:@44155.4]
  input         io_RID, // @[:@44155.4]
  input  [31:0] io_RDATA, // @[:@44155.4]
  input  [1:0]  io_RRESP, // @[:@44155.4]
  input         io_RLAST, // @[:@44155.4]
  input         io_RVALID, // @[:@44155.4]
  output        io_RREADY, // @[:@44155.4]
  output        io_AWID, // @[:@44155.4]
  output [30:0] io_AWADDR, // @[:@44155.4]
  output [7:0]  io_AWLEN, // @[:@44155.4]
  output [2:0]  io_AWSIZE, // @[:@44155.4]
  output [1:0]  io_AWBURST, // @[:@44155.4]
  output        io_AWLOCK, // @[:@44155.4]
  output [3:0]  io_AWCACHE, // @[:@44155.4]
  output [2:0]  io_AWPROT, // @[:@44155.4]
  output [3:0]  io_AWQOS, // @[:@44155.4]
  output [3:0]  io_AWREGION, // @[:@44155.4]
  output        io_AWVALID, // @[:@44155.4]
  input         io_AWREADY, // @[:@44155.4]
  output        io_WID, // @[:@44155.4]
  output [31:0] io_WDATA, // @[:@44155.4]
  output [3:0]  io_WSTRB, // @[:@44155.4]
  output        io_WLAST, // @[:@44155.4]
  output        io_WVALID, // @[:@44155.4]
  input         io_WREADY, // @[:@44155.4]
  input         io_BID, // @[:@44155.4]
  input  [1:0]  io_BRESP, // @[:@44155.4]
  input         io_BVALID, // @[:@44155.4]
  output        io_BREADY, // @[:@44155.4]
  input         io_bbStartSignals_0, // @[:@44155.4]
  input         io_bbStartSignals_1, // @[:@44155.4]
  output        io_bbReadyToPrevious_0, // @[:@44155.4]
  output        io_bbReadyToPrevious_1, // @[:@44155.4]
  output        io_previousAndLoadPorts_0_ready, // @[:@44155.4]
  input         io_previousAndLoadPorts_0_valid, // @[:@44155.4]
  input  [30:0] io_previousAndLoadPorts_0_bits, // @[:@44155.4]
  input         io_nextAndLoadPorts_0_ready, // @[:@44155.4]
  output        io_nextAndLoadPorts_0_valid, // @[:@44155.4]
  output [31:0] io_nextAndLoadPorts_0_bits, // @[:@44155.4]
  output        io_previousAndStoreAddressPorts_0_ready, // @[:@44155.4]
  input         io_previousAndStoreAddressPorts_0_valid, // @[:@44155.4]
  input  [30:0] io_previousAndStoreAddressPorts_0_bits, // @[:@44155.4]
  output        io_previousAndStoreDataPorts_0_ready, // @[:@44155.4]
  input         io_previousAndStoreDataPorts_0_valid, // @[:@44155.4]
  input  [31:0] io_previousAndStoreDataPorts_0_bits, // @[:@44155.4]
  output        io_queueIsEmpty // @[:@44155.4]
);
  wire  storeQ_clock; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_reset; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_bbStart; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_bbStoreOffsets_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_bbNumStores; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_storeTail; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_storeHead; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeEmpty; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_loadTail; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_loadHead; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadEmpty; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadAddressDone_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_loadDataDone_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_loadAddressQueue_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrDone_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataDone_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrQueue_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_1; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_2; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_3; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_4; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_5; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_6; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_7; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_8; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_9; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_10; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_11; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_12; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_13; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_14; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataQueue_15; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeDataEnable_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_dataFromStorePorts_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeAddrEnable_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_addressFromStorePorts_0; // @[LSQAXI.scala 130:22:@44196.4]
  wire [30:0] storeQ_io_storeAddrToMem; // @[LSQAXI.scala 130:22:@44196.4]
  wire [31:0] storeQ_io_storeDataToMem; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeQIdxOut_ready; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeQIdxOut_valid; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_storeQIdxOut_bits; // @[LSQAXI.scala 130:22:@44196.4]
  wire [3:0] storeQ_io_storeQIdxIn; // @[LSQAXI.scala 130:22:@44196.4]
  wire  storeQ_io_storeQIdxInValid; // @[LSQAXI.scala 130:22:@44196.4]
  wire  loadQ_clock; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_reset; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_bbStart; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_bbLoadOffsets_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_bbNumLoads; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_loadTail; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_loadHead; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadEmpty; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_storeTail; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_storeHead; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeEmpty; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeAddrDone_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_storeDataDone_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_storeAddrQueue_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_storeDataQueue_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrDone_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadDataDone_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_1; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_2; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_3; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_4; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_5; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_6; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_7; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_8; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_9; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_10; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_11; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_12; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_13; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_14; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrQueue_15; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadAddrEnable_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_addrFromLoadPorts_0; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadPorts_0_ready; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadPorts_0_valid; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_loadPorts_0_bits; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_loadDataFromMem; // @[LSQAXI.scala 131:21:@44199.4]
  wire [30:0] loadQ_io_loadAddrToMem; // @[LSQAXI.scala 131:21:@44199.4]
  wire [31:0] loadQ_io_loadQIdxForDataIn; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadQIdxForDataInValid; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadQIdxForAddrOut_ready; // @[LSQAXI.scala 131:21:@44199.4]
  wire  loadQ_io_loadQIdxForAddrOut_valid; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] loadQ_io_loadQIdxForAddrOut_bits; // @[LSQAXI.scala 131:21:@44199.4]
  wire [3:0] GA_io_bbLoadOffsets_0; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_1; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_2; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_3; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_4; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_5; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_6; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_7; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_8; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_9; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_10; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_11; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_12; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_13; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_14; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbLoadOffsets_15; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_bbNumLoads; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_loadTail; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_loadHead; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_loadEmpty; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_0; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_1; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_2; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_3; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_4; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_5; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_6; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_7; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_8; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_9; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_10; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_11; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_12; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_13; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_14; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_bbStoreOffsets_15; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_bbNumStores; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_storeTail; // @[LSQAXI.scala 132:18:@44202.4]
  wire [3:0] GA_io_storeHead; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_storeEmpty; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_bbStart; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_bbStartSignals_0; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_bbStartSignals_1; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_readyToPrevious_0; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_readyToPrevious_1; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_loadPortsEnable_0; // @[LSQAXI.scala 132:18:@44202.4]
  wire  GA_io_storePortsEnable_0; // @[LSQAXI.scala 132:18:@44202.4]
  wire  AXIWr_clock; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_reset; // @[LSQAXI.scala 133:21:@44205.4]
  wire [30:0] AXIWr_io_storeAddrToMem; // @[LSQAXI.scala 133:21:@44205.4]
  wire [31:0] AXIWr_io_storeDataToMem; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_storeQIdxInToAW_ready; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_storeQIdxInToAW_valid; // @[LSQAXI.scala 133:21:@44205.4]
  wire [3:0] AXIWr_io_storeQIdxInToAW_bits; // @[LSQAXI.scala 133:21:@44205.4]
  wire [3:0] AXIWr_io_storeQIdxOutFromAW; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_storeQIdxOutFromAWValid; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_AWID; // @[LSQAXI.scala 133:21:@44205.4]
  wire [30:0] AXIWr_io_AWADDR; // @[LSQAXI.scala 133:21:@44205.4]
  wire [7:0] AXIWr_io_AWLEN; // @[LSQAXI.scala 133:21:@44205.4]
  wire [2:0] AXIWr_io_AWSIZE; // @[LSQAXI.scala 133:21:@44205.4]
  wire [1:0] AXIWr_io_AWBURST; // @[LSQAXI.scala 133:21:@44205.4]
  wire [2:0] AXIWr_io_AWPROT; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_AWVALID; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_AWREADY; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_AWLOCK; // @[LSQAXI.scala 133:21:@44205.4]
  wire [3:0] AXIWr_io_AWCACHE; // @[LSQAXI.scala 133:21:@44205.4]
  wire [3:0] AXIWr_io_AWQOS; // @[LSQAXI.scala 133:21:@44205.4]
  wire [3:0] AXIWr_io_AWREGION; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_WID; // @[LSQAXI.scala 133:21:@44205.4]
  wire [31:0] AXIWr_io_WDATA; // @[LSQAXI.scala 133:21:@44205.4]
  wire [3:0] AXIWr_io_WSTRB; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_WLAST; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_WVALID; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_WREADY; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_BID; // @[LSQAXI.scala 133:21:@44205.4]
  wire [1:0] AXIWr_io_BRESP; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_BVALID; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIWr_io_BREADY; // @[LSQAXI.scala 133:21:@44205.4]
  wire  AXIRd_clock; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_reset; // @[LSQAXI.scala 134:21:@44208.4]
  wire [31:0] AXIRd_io_loadDataFromMem; // @[LSQAXI.scala 134:21:@44208.4]
  wire [30:0] AXIRd_io_loadAddrToMem; // @[LSQAXI.scala 134:21:@44208.4]
  wire [31:0] AXIRd_io_loadQIdxForDataOut; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_loadQIdxForDataOutValid; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_loadQIdxForAddrIn_ready; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_loadQIdxForAddrIn_valid; // @[LSQAXI.scala 134:21:@44208.4]
  wire [30:0] AXIRd_io_loadQIdxForAddrIn_bits; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_ARID; // @[LSQAXI.scala 134:21:@44208.4]
  wire [30:0] AXIRd_io_ARADDR; // @[LSQAXI.scala 134:21:@44208.4]
  wire [7:0] AXIRd_io_ARLEN; // @[LSQAXI.scala 134:21:@44208.4]
  wire [2:0] AXIRd_io_ARSIZE; // @[LSQAXI.scala 134:21:@44208.4]
  wire [1:0] AXIRd_io_ARBURST; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_ARLOCK; // @[LSQAXI.scala 134:21:@44208.4]
  wire [3:0] AXIRd_io_ARCACHE; // @[LSQAXI.scala 134:21:@44208.4]
  wire [3:0] AXIRd_io_ARQOS; // @[LSQAXI.scala 134:21:@44208.4]
  wire [3:0] AXIRd_io_ARREGION; // @[LSQAXI.scala 134:21:@44208.4]
  wire [2:0] AXIRd_io_ARPROT; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_ARVALID; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_ARREADY; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_RID; // @[LSQAXI.scala 134:21:@44208.4]
  wire [31:0] AXIRd_io_RDATA; // @[LSQAXI.scala 134:21:@44208.4]
  wire [1:0] AXIRd_io_RRESP; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_RLAST; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_RVALID; // @[LSQAXI.scala 134:21:@44208.4]
  wire  AXIRd_io_RREADY; // @[LSQAXI.scala 134:21:@44208.4]
  wire  LOAD_PORT_LSQ_a_clock; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_reset; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_addrFromPrev_ready; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_addrFromPrev_valid; // @[LSQAXI.scala 138:11:@44211.4]
  wire [30:0] LOAD_PORT_LSQ_a_io_addrFromPrev_bits; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_portEnable; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_dataToNext_ready; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_dataToNext_valid; // @[LSQAXI.scala 138:11:@44211.4]
  wire [31:0] LOAD_PORT_LSQ_a_io_dataToNext_bits; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_loadAddrEnable; // @[LSQAXI.scala 138:11:@44211.4]
  wire [30:0] LOAD_PORT_LSQ_a_io_addrToLoadQueue; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_dataFromLoadQueue_ready; // @[LSQAXI.scala 138:11:@44211.4]
  wire  LOAD_PORT_LSQ_a_io_dataFromLoadQueue_valid; // @[LSQAXI.scala 138:11:@44211.4]
  wire [31:0] LOAD_PORT_LSQ_a_io_dataFromLoadQueue_bits; // @[LSQAXI.scala 138:11:@44211.4]
  wire  STORE_DATA_PORT_LSQ_a_clock; // @[LSQAXI.scala 142:11:@44227.4]
  wire  STORE_DATA_PORT_LSQ_a_reset; // @[LSQAXI.scala 142:11:@44227.4]
  wire  STORE_DATA_PORT_LSQ_a_io_dataFromPrev_ready; // @[LSQAXI.scala 142:11:@44227.4]
  wire  STORE_DATA_PORT_LSQ_a_io_dataFromPrev_valid; // @[LSQAXI.scala 142:11:@44227.4]
  wire [31:0] STORE_DATA_PORT_LSQ_a_io_dataFromPrev_bits; // @[LSQAXI.scala 142:11:@44227.4]
  wire  STORE_DATA_PORT_LSQ_a_io_portEnable; // @[LSQAXI.scala 142:11:@44227.4]
  wire  STORE_DATA_PORT_LSQ_a_io_storeDataEnable; // @[LSQAXI.scala 142:11:@44227.4]
  wire [31:0] STORE_DATA_PORT_LSQ_a_io_dataToStoreQueue; // @[LSQAXI.scala 142:11:@44227.4]
  wire  STORE_ADDR_PORT_LSQ_a_clock; // @[LSQAXI.scala 146:11:@44237.4]
  wire  STORE_ADDR_PORT_LSQ_a_reset; // @[LSQAXI.scala 146:11:@44237.4]
  wire  STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_ready; // @[LSQAXI.scala 146:11:@44237.4]
  wire  STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_valid; // @[LSQAXI.scala 146:11:@44237.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_bits; // @[LSQAXI.scala 146:11:@44237.4]
  wire  STORE_ADDR_PORT_LSQ_a_io_portEnable; // @[LSQAXI.scala 146:11:@44237.4]
  wire  STORE_ADDR_PORT_LSQ_a_io_storeDataEnable; // @[LSQAXI.scala 146:11:@44237.4]
  wire [31:0] STORE_ADDR_PORT_LSQ_a_io_dataToStoreQueue; // @[LSQAXI.scala 146:11:@44237.4]
  wire  storeEmpty; // @[LSQAXI.scala 89:24:@44162.4 LSQAXI.scala 216:14:@44579.4]
  wire  loadEmpty; // @[LSQAXI.scala 95:23:@44168.4 LSQAXI.scala 184:13:@44431.4]
  wire [15:0] storeTail; // @[LSQAXI.scala 87:23:@44160.4 LSQAXI.scala 214:13:@44577.4]
  wire [15:0] storeHead; // @[LSQAXI.scala 88:23:@44161.4 LSQAXI.scala 215:13:@44578.4]
  wire [15:0] loadTail; // @[LSQAXI.scala 93:22:@44166.4 LSQAXI.scala 182:12:@44429.4]
  wire [15:0] loadHead; // @[LSQAXI.scala 94:22:@44167.4 LSQAXI.scala 183:12:@44430.4]
  wire [31:0] sAddressPorts_0_addrToStoreQueue; // @[LSQAXI.scala 145:30:@44240.4 LSQAXI.scala 145:30:@44241.4]
  STORE_QUEUE storeQ ( // @[LSQAXI.scala 130:22:@44196.4]
    .clock(storeQ_clock),
    .reset(storeQ_reset),
    .io_bbStart(storeQ_io_bbStart),
    .io_bbStoreOffsets_0(storeQ_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(storeQ_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(storeQ_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(storeQ_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(storeQ_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(storeQ_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(storeQ_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(storeQ_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(storeQ_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(storeQ_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(storeQ_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(storeQ_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(storeQ_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(storeQ_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(storeQ_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(storeQ_io_bbStoreOffsets_15),
    .io_bbNumStores(storeQ_io_bbNumStores),
    .io_storeTail(storeQ_io_storeTail),
    .io_storeHead(storeQ_io_storeHead),
    .io_storeEmpty(storeQ_io_storeEmpty),
    .io_loadTail(storeQ_io_loadTail),
    .io_loadHead(storeQ_io_loadHead),
    .io_loadEmpty(storeQ_io_loadEmpty),
    .io_loadAddressDone_0(storeQ_io_loadAddressDone_0),
    .io_loadAddressDone_1(storeQ_io_loadAddressDone_1),
    .io_loadAddressDone_2(storeQ_io_loadAddressDone_2),
    .io_loadAddressDone_3(storeQ_io_loadAddressDone_3),
    .io_loadAddressDone_4(storeQ_io_loadAddressDone_4),
    .io_loadAddressDone_5(storeQ_io_loadAddressDone_5),
    .io_loadAddressDone_6(storeQ_io_loadAddressDone_6),
    .io_loadAddressDone_7(storeQ_io_loadAddressDone_7),
    .io_loadAddressDone_8(storeQ_io_loadAddressDone_8),
    .io_loadAddressDone_9(storeQ_io_loadAddressDone_9),
    .io_loadAddressDone_10(storeQ_io_loadAddressDone_10),
    .io_loadAddressDone_11(storeQ_io_loadAddressDone_11),
    .io_loadAddressDone_12(storeQ_io_loadAddressDone_12),
    .io_loadAddressDone_13(storeQ_io_loadAddressDone_13),
    .io_loadAddressDone_14(storeQ_io_loadAddressDone_14),
    .io_loadAddressDone_15(storeQ_io_loadAddressDone_15),
    .io_loadDataDone_0(storeQ_io_loadDataDone_0),
    .io_loadDataDone_1(storeQ_io_loadDataDone_1),
    .io_loadDataDone_2(storeQ_io_loadDataDone_2),
    .io_loadDataDone_3(storeQ_io_loadDataDone_3),
    .io_loadDataDone_4(storeQ_io_loadDataDone_4),
    .io_loadDataDone_5(storeQ_io_loadDataDone_5),
    .io_loadDataDone_6(storeQ_io_loadDataDone_6),
    .io_loadDataDone_7(storeQ_io_loadDataDone_7),
    .io_loadDataDone_8(storeQ_io_loadDataDone_8),
    .io_loadDataDone_9(storeQ_io_loadDataDone_9),
    .io_loadDataDone_10(storeQ_io_loadDataDone_10),
    .io_loadDataDone_11(storeQ_io_loadDataDone_11),
    .io_loadDataDone_12(storeQ_io_loadDataDone_12),
    .io_loadDataDone_13(storeQ_io_loadDataDone_13),
    .io_loadDataDone_14(storeQ_io_loadDataDone_14),
    .io_loadDataDone_15(storeQ_io_loadDataDone_15),
    .io_loadAddressQueue_0(storeQ_io_loadAddressQueue_0),
    .io_loadAddressQueue_1(storeQ_io_loadAddressQueue_1),
    .io_loadAddressQueue_2(storeQ_io_loadAddressQueue_2),
    .io_loadAddressQueue_3(storeQ_io_loadAddressQueue_3),
    .io_loadAddressQueue_4(storeQ_io_loadAddressQueue_4),
    .io_loadAddressQueue_5(storeQ_io_loadAddressQueue_5),
    .io_loadAddressQueue_6(storeQ_io_loadAddressQueue_6),
    .io_loadAddressQueue_7(storeQ_io_loadAddressQueue_7),
    .io_loadAddressQueue_8(storeQ_io_loadAddressQueue_8),
    .io_loadAddressQueue_9(storeQ_io_loadAddressQueue_9),
    .io_loadAddressQueue_10(storeQ_io_loadAddressQueue_10),
    .io_loadAddressQueue_11(storeQ_io_loadAddressQueue_11),
    .io_loadAddressQueue_12(storeQ_io_loadAddressQueue_12),
    .io_loadAddressQueue_13(storeQ_io_loadAddressQueue_13),
    .io_loadAddressQueue_14(storeQ_io_loadAddressQueue_14),
    .io_loadAddressQueue_15(storeQ_io_loadAddressQueue_15),
    .io_storeAddrDone_0(storeQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(storeQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(storeQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(storeQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(storeQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(storeQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(storeQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(storeQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(storeQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(storeQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(storeQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(storeQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(storeQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(storeQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(storeQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(storeQ_io_storeAddrDone_15),
    .io_storeDataDone_0(storeQ_io_storeDataDone_0),
    .io_storeDataDone_1(storeQ_io_storeDataDone_1),
    .io_storeDataDone_2(storeQ_io_storeDataDone_2),
    .io_storeDataDone_3(storeQ_io_storeDataDone_3),
    .io_storeDataDone_4(storeQ_io_storeDataDone_4),
    .io_storeDataDone_5(storeQ_io_storeDataDone_5),
    .io_storeDataDone_6(storeQ_io_storeDataDone_6),
    .io_storeDataDone_7(storeQ_io_storeDataDone_7),
    .io_storeDataDone_8(storeQ_io_storeDataDone_8),
    .io_storeDataDone_9(storeQ_io_storeDataDone_9),
    .io_storeDataDone_10(storeQ_io_storeDataDone_10),
    .io_storeDataDone_11(storeQ_io_storeDataDone_11),
    .io_storeDataDone_12(storeQ_io_storeDataDone_12),
    .io_storeDataDone_13(storeQ_io_storeDataDone_13),
    .io_storeDataDone_14(storeQ_io_storeDataDone_14),
    .io_storeDataDone_15(storeQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(storeQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(storeQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(storeQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(storeQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(storeQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(storeQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(storeQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(storeQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(storeQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(storeQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(storeQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(storeQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(storeQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(storeQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(storeQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(storeQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(storeQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(storeQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(storeQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(storeQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(storeQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(storeQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(storeQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(storeQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(storeQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(storeQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(storeQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(storeQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(storeQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(storeQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(storeQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(storeQ_io_storeDataQueue_15),
    .io_storeDataEnable_0(storeQ_io_storeDataEnable_0),
    .io_dataFromStorePorts_0(storeQ_io_dataFromStorePorts_0),
    .io_storeAddrEnable_0(storeQ_io_storeAddrEnable_0),
    .io_addressFromStorePorts_0(storeQ_io_addressFromStorePorts_0),
    .io_storeAddrToMem(storeQ_io_storeAddrToMem),
    .io_storeDataToMem(storeQ_io_storeDataToMem),
    .io_storeQIdxOut_ready(storeQ_io_storeQIdxOut_ready),
    .io_storeQIdxOut_valid(storeQ_io_storeQIdxOut_valid),
    .io_storeQIdxOut_bits(storeQ_io_storeQIdxOut_bits),
    .io_storeQIdxIn(storeQ_io_storeQIdxIn),
    .io_storeQIdxInValid(storeQ_io_storeQIdxInValid)
  );
  LOAD_QUEUE loadQ ( // @[LSQAXI.scala 131:21:@44199.4]
    .clock(loadQ_clock),
    .reset(loadQ_reset),
    .io_bbStart(loadQ_io_bbStart),
    .io_bbLoadOffsets_0(loadQ_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(loadQ_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(loadQ_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(loadQ_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(loadQ_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(loadQ_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(loadQ_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(loadQ_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(loadQ_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(loadQ_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(loadQ_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(loadQ_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(loadQ_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(loadQ_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(loadQ_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(loadQ_io_bbLoadOffsets_15),
    .io_bbNumLoads(loadQ_io_bbNumLoads),
    .io_loadTail(loadQ_io_loadTail),
    .io_loadHead(loadQ_io_loadHead),
    .io_loadEmpty(loadQ_io_loadEmpty),
    .io_storeTail(loadQ_io_storeTail),
    .io_storeHead(loadQ_io_storeHead),
    .io_storeEmpty(loadQ_io_storeEmpty),
    .io_storeAddrDone_0(loadQ_io_storeAddrDone_0),
    .io_storeAddrDone_1(loadQ_io_storeAddrDone_1),
    .io_storeAddrDone_2(loadQ_io_storeAddrDone_2),
    .io_storeAddrDone_3(loadQ_io_storeAddrDone_3),
    .io_storeAddrDone_4(loadQ_io_storeAddrDone_4),
    .io_storeAddrDone_5(loadQ_io_storeAddrDone_5),
    .io_storeAddrDone_6(loadQ_io_storeAddrDone_6),
    .io_storeAddrDone_7(loadQ_io_storeAddrDone_7),
    .io_storeAddrDone_8(loadQ_io_storeAddrDone_8),
    .io_storeAddrDone_9(loadQ_io_storeAddrDone_9),
    .io_storeAddrDone_10(loadQ_io_storeAddrDone_10),
    .io_storeAddrDone_11(loadQ_io_storeAddrDone_11),
    .io_storeAddrDone_12(loadQ_io_storeAddrDone_12),
    .io_storeAddrDone_13(loadQ_io_storeAddrDone_13),
    .io_storeAddrDone_14(loadQ_io_storeAddrDone_14),
    .io_storeAddrDone_15(loadQ_io_storeAddrDone_15),
    .io_storeDataDone_0(loadQ_io_storeDataDone_0),
    .io_storeDataDone_1(loadQ_io_storeDataDone_1),
    .io_storeDataDone_2(loadQ_io_storeDataDone_2),
    .io_storeDataDone_3(loadQ_io_storeDataDone_3),
    .io_storeDataDone_4(loadQ_io_storeDataDone_4),
    .io_storeDataDone_5(loadQ_io_storeDataDone_5),
    .io_storeDataDone_6(loadQ_io_storeDataDone_6),
    .io_storeDataDone_7(loadQ_io_storeDataDone_7),
    .io_storeDataDone_8(loadQ_io_storeDataDone_8),
    .io_storeDataDone_9(loadQ_io_storeDataDone_9),
    .io_storeDataDone_10(loadQ_io_storeDataDone_10),
    .io_storeDataDone_11(loadQ_io_storeDataDone_11),
    .io_storeDataDone_12(loadQ_io_storeDataDone_12),
    .io_storeDataDone_13(loadQ_io_storeDataDone_13),
    .io_storeDataDone_14(loadQ_io_storeDataDone_14),
    .io_storeDataDone_15(loadQ_io_storeDataDone_15),
    .io_storeAddrQueue_0(loadQ_io_storeAddrQueue_0),
    .io_storeAddrQueue_1(loadQ_io_storeAddrQueue_1),
    .io_storeAddrQueue_2(loadQ_io_storeAddrQueue_2),
    .io_storeAddrQueue_3(loadQ_io_storeAddrQueue_3),
    .io_storeAddrQueue_4(loadQ_io_storeAddrQueue_4),
    .io_storeAddrQueue_5(loadQ_io_storeAddrQueue_5),
    .io_storeAddrQueue_6(loadQ_io_storeAddrQueue_6),
    .io_storeAddrQueue_7(loadQ_io_storeAddrQueue_7),
    .io_storeAddrQueue_8(loadQ_io_storeAddrQueue_8),
    .io_storeAddrQueue_9(loadQ_io_storeAddrQueue_9),
    .io_storeAddrQueue_10(loadQ_io_storeAddrQueue_10),
    .io_storeAddrQueue_11(loadQ_io_storeAddrQueue_11),
    .io_storeAddrQueue_12(loadQ_io_storeAddrQueue_12),
    .io_storeAddrQueue_13(loadQ_io_storeAddrQueue_13),
    .io_storeAddrQueue_14(loadQ_io_storeAddrQueue_14),
    .io_storeAddrQueue_15(loadQ_io_storeAddrQueue_15),
    .io_storeDataQueue_0(loadQ_io_storeDataQueue_0),
    .io_storeDataQueue_1(loadQ_io_storeDataQueue_1),
    .io_storeDataQueue_2(loadQ_io_storeDataQueue_2),
    .io_storeDataQueue_3(loadQ_io_storeDataQueue_3),
    .io_storeDataQueue_4(loadQ_io_storeDataQueue_4),
    .io_storeDataQueue_5(loadQ_io_storeDataQueue_5),
    .io_storeDataQueue_6(loadQ_io_storeDataQueue_6),
    .io_storeDataQueue_7(loadQ_io_storeDataQueue_7),
    .io_storeDataQueue_8(loadQ_io_storeDataQueue_8),
    .io_storeDataQueue_9(loadQ_io_storeDataQueue_9),
    .io_storeDataQueue_10(loadQ_io_storeDataQueue_10),
    .io_storeDataQueue_11(loadQ_io_storeDataQueue_11),
    .io_storeDataQueue_12(loadQ_io_storeDataQueue_12),
    .io_storeDataQueue_13(loadQ_io_storeDataQueue_13),
    .io_storeDataQueue_14(loadQ_io_storeDataQueue_14),
    .io_storeDataQueue_15(loadQ_io_storeDataQueue_15),
    .io_loadAddrDone_0(loadQ_io_loadAddrDone_0),
    .io_loadAddrDone_1(loadQ_io_loadAddrDone_1),
    .io_loadAddrDone_2(loadQ_io_loadAddrDone_2),
    .io_loadAddrDone_3(loadQ_io_loadAddrDone_3),
    .io_loadAddrDone_4(loadQ_io_loadAddrDone_4),
    .io_loadAddrDone_5(loadQ_io_loadAddrDone_5),
    .io_loadAddrDone_6(loadQ_io_loadAddrDone_6),
    .io_loadAddrDone_7(loadQ_io_loadAddrDone_7),
    .io_loadAddrDone_8(loadQ_io_loadAddrDone_8),
    .io_loadAddrDone_9(loadQ_io_loadAddrDone_9),
    .io_loadAddrDone_10(loadQ_io_loadAddrDone_10),
    .io_loadAddrDone_11(loadQ_io_loadAddrDone_11),
    .io_loadAddrDone_12(loadQ_io_loadAddrDone_12),
    .io_loadAddrDone_13(loadQ_io_loadAddrDone_13),
    .io_loadAddrDone_14(loadQ_io_loadAddrDone_14),
    .io_loadAddrDone_15(loadQ_io_loadAddrDone_15),
    .io_loadDataDone_0(loadQ_io_loadDataDone_0),
    .io_loadDataDone_1(loadQ_io_loadDataDone_1),
    .io_loadDataDone_2(loadQ_io_loadDataDone_2),
    .io_loadDataDone_3(loadQ_io_loadDataDone_3),
    .io_loadDataDone_4(loadQ_io_loadDataDone_4),
    .io_loadDataDone_5(loadQ_io_loadDataDone_5),
    .io_loadDataDone_6(loadQ_io_loadDataDone_6),
    .io_loadDataDone_7(loadQ_io_loadDataDone_7),
    .io_loadDataDone_8(loadQ_io_loadDataDone_8),
    .io_loadDataDone_9(loadQ_io_loadDataDone_9),
    .io_loadDataDone_10(loadQ_io_loadDataDone_10),
    .io_loadDataDone_11(loadQ_io_loadDataDone_11),
    .io_loadDataDone_12(loadQ_io_loadDataDone_12),
    .io_loadDataDone_13(loadQ_io_loadDataDone_13),
    .io_loadDataDone_14(loadQ_io_loadDataDone_14),
    .io_loadDataDone_15(loadQ_io_loadDataDone_15),
    .io_loadAddrQueue_0(loadQ_io_loadAddrQueue_0),
    .io_loadAddrQueue_1(loadQ_io_loadAddrQueue_1),
    .io_loadAddrQueue_2(loadQ_io_loadAddrQueue_2),
    .io_loadAddrQueue_3(loadQ_io_loadAddrQueue_3),
    .io_loadAddrQueue_4(loadQ_io_loadAddrQueue_4),
    .io_loadAddrQueue_5(loadQ_io_loadAddrQueue_5),
    .io_loadAddrQueue_6(loadQ_io_loadAddrQueue_6),
    .io_loadAddrQueue_7(loadQ_io_loadAddrQueue_7),
    .io_loadAddrQueue_8(loadQ_io_loadAddrQueue_8),
    .io_loadAddrQueue_9(loadQ_io_loadAddrQueue_9),
    .io_loadAddrQueue_10(loadQ_io_loadAddrQueue_10),
    .io_loadAddrQueue_11(loadQ_io_loadAddrQueue_11),
    .io_loadAddrQueue_12(loadQ_io_loadAddrQueue_12),
    .io_loadAddrQueue_13(loadQ_io_loadAddrQueue_13),
    .io_loadAddrQueue_14(loadQ_io_loadAddrQueue_14),
    .io_loadAddrQueue_15(loadQ_io_loadAddrQueue_15),
    .io_loadAddrEnable_0(loadQ_io_loadAddrEnable_0),
    .io_addrFromLoadPorts_0(loadQ_io_addrFromLoadPorts_0),
    .io_loadPorts_0_ready(loadQ_io_loadPorts_0_ready),
    .io_loadPorts_0_valid(loadQ_io_loadPorts_0_valid),
    .io_loadPorts_0_bits(loadQ_io_loadPorts_0_bits),
    .io_loadDataFromMem(loadQ_io_loadDataFromMem),
    .io_loadAddrToMem(loadQ_io_loadAddrToMem),
    .io_loadQIdxForDataIn(loadQ_io_loadQIdxForDataIn),
    .io_loadQIdxForDataInValid(loadQ_io_loadQIdxForDataInValid),
    .io_loadQIdxForAddrOut_ready(loadQ_io_loadQIdxForAddrOut_ready),
    .io_loadQIdxForAddrOut_valid(loadQ_io_loadQIdxForAddrOut_valid),
    .io_loadQIdxForAddrOut_bits(loadQ_io_loadQIdxForAddrOut_bits)
  );
  GROUP_ALLOCATOR_LSQ_a GA ( // @[LSQAXI.scala 132:18:@44202.4]
    .io_bbLoadOffsets_0(GA_io_bbLoadOffsets_0),
    .io_bbLoadOffsets_1(GA_io_bbLoadOffsets_1),
    .io_bbLoadOffsets_2(GA_io_bbLoadOffsets_2),
    .io_bbLoadOffsets_3(GA_io_bbLoadOffsets_3),
    .io_bbLoadOffsets_4(GA_io_bbLoadOffsets_4),
    .io_bbLoadOffsets_5(GA_io_bbLoadOffsets_5),
    .io_bbLoadOffsets_6(GA_io_bbLoadOffsets_6),
    .io_bbLoadOffsets_7(GA_io_bbLoadOffsets_7),
    .io_bbLoadOffsets_8(GA_io_bbLoadOffsets_8),
    .io_bbLoadOffsets_9(GA_io_bbLoadOffsets_9),
    .io_bbLoadOffsets_10(GA_io_bbLoadOffsets_10),
    .io_bbLoadOffsets_11(GA_io_bbLoadOffsets_11),
    .io_bbLoadOffsets_12(GA_io_bbLoadOffsets_12),
    .io_bbLoadOffsets_13(GA_io_bbLoadOffsets_13),
    .io_bbLoadOffsets_14(GA_io_bbLoadOffsets_14),
    .io_bbLoadOffsets_15(GA_io_bbLoadOffsets_15),
    .io_bbNumLoads(GA_io_bbNumLoads),
    .io_loadTail(GA_io_loadTail),
    .io_loadHead(GA_io_loadHead),
    .io_loadEmpty(GA_io_loadEmpty),
    .io_bbStoreOffsets_0(GA_io_bbStoreOffsets_0),
    .io_bbStoreOffsets_1(GA_io_bbStoreOffsets_1),
    .io_bbStoreOffsets_2(GA_io_bbStoreOffsets_2),
    .io_bbStoreOffsets_3(GA_io_bbStoreOffsets_3),
    .io_bbStoreOffsets_4(GA_io_bbStoreOffsets_4),
    .io_bbStoreOffsets_5(GA_io_bbStoreOffsets_5),
    .io_bbStoreOffsets_6(GA_io_bbStoreOffsets_6),
    .io_bbStoreOffsets_7(GA_io_bbStoreOffsets_7),
    .io_bbStoreOffsets_8(GA_io_bbStoreOffsets_8),
    .io_bbStoreOffsets_9(GA_io_bbStoreOffsets_9),
    .io_bbStoreOffsets_10(GA_io_bbStoreOffsets_10),
    .io_bbStoreOffsets_11(GA_io_bbStoreOffsets_11),
    .io_bbStoreOffsets_12(GA_io_bbStoreOffsets_12),
    .io_bbStoreOffsets_13(GA_io_bbStoreOffsets_13),
    .io_bbStoreOffsets_14(GA_io_bbStoreOffsets_14),
    .io_bbStoreOffsets_15(GA_io_bbStoreOffsets_15),
    .io_bbNumStores(GA_io_bbNumStores),
    .io_storeTail(GA_io_storeTail),
    .io_storeHead(GA_io_storeHead),
    .io_storeEmpty(GA_io_storeEmpty),
    .io_bbStart(GA_io_bbStart),
    .io_bbStartSignals_0(GA_io_bbStartSignals_0),
    .io_bbStartSignals_1(GA_io_bbStartSignals_1),
    .io_readyToPrevious_0(GA_io_readyToPrevious_0),
    .io_readyToPrevious_1(GA_io_readyToPrevious_1),
    .io_loadPortsEnable_0(GA_io_loadPortsEnable_0),
    .io_storePortsEnable_0(GA_io_storePortsEnable_0)
  );
  AXI_WRITE AXIWr ( // @[LSQAXI.scala 133:21:@44205.4]
    .clock(AXIWr_clock),
    .reset(AXIWr_reset),
    .io_storeAddrToMem(AXIWr_io_storeAddrToMem),
    .io_storeDataToMem(AXIWr_io_storeDataToMem),
    .io_storeQIdxInToAW_ready(AXIWr_io_storeQIdxInToAW_ready),
    .io_storeQIdxInToAW_valid(AXIWr_io_storeQIdxInToAW_valid),
    .io_storeQIdxInToAW_bits(AXIWr_io_storeQIdxInToAW_bits),
    .io_storeQIdxOutFromAW(AXIWr_io_storeQIdxOutFromAW),
    .io_storeQIdxOutFromAWValid(AXIWr_io_storeQIdxOutFromAWValid),
    .io_AWID(AXIWr_io_AWID),
    .io_AWADDR(AXIWr_io_AWADDR),
    .io_AWLEN(AXIWr_io_AWLEN),
    .io_AWSIZE(AXIWr_io_AWSIZE),
    .io_AWBURST(AXIWr_io_AWBURST),
    .io_AWPROT(AXIWr_io_AWPROT),
    .io_AWVALID(AXIWr_io_AWVALID),
    .io_AWREADY(AXIWr_io_AWREADY),
    .io_AWLOCK(AXIWr_io_AWLOCK),
    .io_AWCACHE(AXIWr_io_AWCACHE),
    .io_AWQOS(AXIWr_io_AWQOS),
    .io_AWREGION(AXIWr_io_AWREGION),
    .io_WID(AXIWr_io_WID),
    .io_WDATA(AXIWr_io_WDATA),
    .io_WSTRB(AXIWr_io_WSTRB),
    .io_WLAST(AXIWr_io_WLAST),
    .io_WVALID(AXIWr_io_WVALID),
    .io_WREADY(AXIWr_io_WREADY),
    .io_BID(AXIWr_io_BID),
    .io_BRESP(AXIWr_io_BRESP),
    .io_BVALID(AXIWr_io_BVALID),
    .io_BREADY(AXIWr_io_BREADY)
  );
  AXI_READ AXIRd ( // @[LSQAXI.scala 134:21:@44208.4]
    .clock(AXIRd_clock),
    .reset(AXIRd_reset),
    .io_loadDataFromMem(AXIRd_io_loadDataFromMem),
    .io_loadAddrToMem(AXIRd_io_loadAddrToMem),
    .io_loadQIdxForDataOut(AXIRd_io_loadQIdxForDataOut),
    .io_loadQIdxForDataOutValid(AXIRd_io_loadQIdxForDataOutValid),
    .io_loadQIdxForAddrIn_ready(AXIRd_io_loadQIdxForAddrIn_ready),
    .io_loadQIdxForAddrIn_valid(AXIRd_io_loadQIdxForAddrIn_valid),
    .io_loadQIdxForAddrIn_bits(AXIRd_io_loadQIdxForAddrIn_bits),
    .io_ARID(AXIRd_io_ARID),
    .io_ARADDR(AXIRd_io_ARADDR),
    .io_ARLEN(AXIRd_io_ARLEN),
    .io_ARSIZE(AXIRd_io_ARSIZE),
    .io_ARBURST(AXIRd_io_ARBURST),
    .io_ARLOCK(AXIRd_io_ARLOCK),
    .io_ARCACHE(AXIRd_io_ARCACHE),
    .io_ARQOS(AXIRd_io_ARQOS),
    .io_ARREGION(AXIRd_io_ARREGION),
    .io_ARPROT(AXIRd_io_ARPROT),
    .io_ARVALID(AXIRd_io_ARVALID),
    .io_ARREADY(AXIRd_io_ARREADY),
    .io_RID(AXIRd_io_RID),
    .io_RDATA(AXIRd_io_RDATA),
    .io_RRESP(AXIRd_io_RRESP),
    .io_RLAST(AXIRd_io_RLAST),
    .io_RVALID(AXIRd_io_RVALID),
    .io_RREADY(AXIRd_io_RREADY)
  );
  LOAD_PORT_LSQ_a LOAD_PORT_LSQ_a ( // @[LSQAXI.scala 138:11:@44211.4]
    .clock(LOAD_PORT_LSQ_a_clock),
    .reset(LOAD_PORT_LSQ_a_reset),
    .io_addrFromPrev_ready(LOAD_PORT_LSQ_a_io_addrFromPrev_ready),
    .io_addrFromPrev_valid(LOAD_PORT_LSQ_a_io_addrFromPrev_valid),
    .io_addrFromPrev_bits(LOAD_PORT_LSQ_a_io_addrFromPrev_bits),
    .io_portEnable(LOAD_PORT_LSQ_a_io_portEnable),
    .io_dataToNext_ready(LOAD_PORT_LSQ_a_io_dataToNext_ready),
    .io_dataToNext_valid(LOAD_PORT_LSQ_a_io_dataToNext_valid),
    .io_dataToNext_bits(LOAD_PORT_LSQ_a_io_dataToNext_bits),
    .io_loadAddrEnable(LOAD_PORT_LSQ_a_io_loadAddrEnable),
    .io_addrToLoadQueue(LOAD_PORT_LSQ_a_io_addrToLoadQueue),
    .io_dataFromLoadQueue_ready(LOAD_PORT_LSQ_a_io_dataFromLoadQueue_ready),
    .io_dataFromLoadQueue_valid(LOAD_PORT_LSQ_a_io_dataFromLoadQueue_valid),
    .io_dataFromLoadQueue_bits(LOAD_PORT_LSQ_a_io_dataFromLoadQueue_bits)
  );
  STORE_DATA_PORT_LSQ_a STORE_DATA_PORT_LSQ_a ( // @[LSQAXI.scala 142:11:@44227.4]
    .clock(STORE_DATA_PORT_LSQ_a_clock),
    .reset(STORE_DATA_PORT_LSQ_a_reset),
    .io_dataFromPrev_ready(STORE_DATA_PORT_LSQ_a_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_DATA_PORT_LSQ_a_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_DATA_PORT_LSQ_a_io_dataFromPrev_bits),
    .io_portEnable(STORE_DATA_PORT_LSQ_a_io_portEnable),
    .io_storeDataEnable(STORE_DATA_PORT_LSQ_a_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_DATA_PORT_LSQ_a_io_dataToStoreQueue)
  );
  STORE_DATA_PORT_LSQ_a STORE_ADDR_PORT_LSQ_a ( // @[LSQAXI.scala 146:11:@44237.4]
    .clock(STORE_ADDR_PORT_LSQ_a_clock),
    .reset(STORE_ADDR_PORT_LSQ_a_reset),
    .io_dataFromPrev_ready(STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_ready),
    .io_dataFromPrev_valid(STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_valid),
    .io_dataFromPrev_bits(STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_bits),
    .io_portEnable(STORE_ADDR_PORT_LSQ_a_io_portEnable),
    .io_storeDataEnable(STORE_ADDR_PORT_LSQ_a_io_storeDataEnable),
    .io_dataToStoreQueue(STORE_ADDR_PORT_LSQ_a_io_dataToStoreQueue)
  );
  assign storeEmpty = storeQ_io_storeEmpty; // @[LSQAXI.scala 89:24:@44162.4 LSQAXI.scala 216:14:@44579.4]
  assign loadEmpty = loadQ_io_loadEmpty; // @[LSQAXI.scala 95:23:@44168.4 LSQAXI.scala 184:13:@44431.4]
  assign storeTail = {{12'd0}, storeQ_io_storeTail}; // @[LSQAXI.scala 87:23:@44160.4 LSQAXI.scala 214:13:@44577.4]
  assign storeHead = {{12'd0}, storeQ_io_storeHead}; // @[LSQAXI.scala 88:23:@44161.4 LSQAXI.scala 215:13:@44578.4]
  assign loadTail = {{12'd0}, loadQ_io_loadTail}; // @[LSQAXI.scala 93:22:@44166.4 LSQAXI.scala 182:12:@44429.4]
  assign loadHead = {{12'd0}, loadQ_io_loadHead}; // @[LSQAXI.scala 94:22:@44167.4 LSQAXI.scala 183:12:@44430.4]
  assign sAddressPorts_0_addrToStoreQueue = STORE_ADDR_PORT_LSQ_a_io_dataToStoreQueue; // @[LSQAXI.scala 145:30:@44240.4 LSQAXI.scala 145:30:@44241.4]
  assign io_ARID = AXIRd_io_ARID; // @[LSQAXI.scala 244:11:@44662.4]
  assign io_ARADDR = AXIRd_io_ARADDR; // @[LSQAXI.scala 245:13:@44663.4]
  assign io_ARLEN = AXIRd_io_ARLEN; // @[LSQAXI.scala 246:12:@44664.4]
  assign io_ARSIZE = AXIRd_io_ARSIZE; // @[LSQAXI.scala 247:13:@44665.4]
  assign io_ARBURST = AXIRd_io_ARBURST; // @[LSQAXI.scala 248:14:@44666.4]
  assign io_ARLOCK = AXIRd_io_ARLOCK; // @[LSQAXI.scala 249:13:@44667.4]
  assign io_ARCACHE = AXIRd_io_ARCACHE; // @[LSQAXI.scala 250:14:@44668.4]
  assign io_ARPROT = AXIRd_io_ARPROT; // @[LSQAXI.scala 251:13:@44669.4]
  assign io_ARQOS = AXIRd_io_ARQOS; // @[LSQAXI.scala 252:12:@44670.4]
  assign io_ARREGION = AXIRd_io_ARREGION; // @[LSQAXI.scala 253:15:@44671.4]
  assign io_ARVALID = AXIRd_io_ARVALID; // @[LSQAXI.scala 254:14:@44672.4]
  assign io_RREADY = AXIRd_io_RREADY; // @[LSQAXI.scala 263:13:@44679.4]
  assign io_AWID = AXIWr_io_AWID; // @[LSQAXI.scala 275:11:@44687.4]
  assign io_AWADDR = AXIWr_io_AWADDR; // @[LSQAXI.scala 276:13:@44688.4]
  assign io_AWLEN = AXIWr_io_AWLEN; // @[LSQAXI.scala 277:12:@44689.4]
  assign io_AWSIZE = AXIWr_io_AWSIZE; // @[LSQAXI.scala 278:13:@44690.4]
  assign io_AWBURST = AXIWr_io_AWBURST; // @[LSQAXI.scala 279:14:@44691.4]
  assign io_AWLOCK = AXIWr_io_AWLOCK; // @[LSQAXI.scala 280:13:@44692.4]
  assign io_AWCACHE = AXIWr_io_AWCACHE; // @[LSQAXI.scala 281:14:@44693.4]
  assign io_AWPROT = AXIWr_io_AWPROT; // @[LSQAXI.scala 282:13:@44694.4]
  assign io_AWQOS = AXIWr_io_AWQOS; // @[LSQAXI.scala 283:12:@44695.4]
  assign io_AWREGION = AXIWr_io_AWREGION; // @[LSQAXI.scala 284:15:@44696.4]
  assign io_AWVALID = AXIWr_io_AWVALID; // @[LSQAXI.scala 285:14:@44697.4]
  assign io_WID = AXIWr_io_WID; // @[LSQAXI.scala 288:10:@44699.4]
  assign io_WDATA = AXIWr_io_WDATA; // @[LSQAXI.scala 289:12:@44700.4]
  assign io_WSTRB = AXIWr_io_WSTRB; // @[LSQAXI.scala 290:12:@44701.4]
  assign io_WLAST = AXIWr_io_WLAST; // @[LSQAXI.scala 291:12:@44702.4]
  assign io_WVALID = AXIWr_io_WVALID; // @[LSQAXI.scala 292:13:@44703.4]
  assign io_BREADY = AXIWr_io_BREADY; // @[LSQAXI.scala 298:13:@44708.4]
  assign io_bbReadyToPrevious_0 = GA_io_readyToPrevious_0; // @[LSQAXI.scala 166:24:@44324.4]
  assign io_bbReadyToPrevious_1 = GA_io_readyToPrevious_1; // @[LSQAXI.scala 166:24:@44325.4]
  assign io_previousAndLoadPorts_0_ready = LOAD_PORT_LSQ_a_io_addrFromPrev_ready; // @[LSQAXI.scala 301:28:@44711.4]
  assign io_nextAndLoadPorts_0_valid = LOAD_PORT_LSQ_a_io_dataToNext_valid; // @[LSQAXI.scala 303:28:@44714.4]
  assign io_nextAndLoadPorts_0_bits = LOAD_PORT_LSQ_a_io_dataToNext_bits; // @[LSQAXI.scala 303:28:@44713.4]
  assign io_previousAndStoreAddressPorts_0_ready = STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_ready; // @[LSQAXI.scala 317:35:@44729.4]
  assign io_previousAndStoreDataPorts_0_ready = STORE_DATA_PORT_LSQ_a_io_dataFromPrev_ready; // @[LSQAXI.scala 312:32:@44723.4]
  assign io_queueIsEmpty = storeEmpty & loadEmpty; // @[LSQAXI.scala 149:19:@44248.4]
  assign storeQ_clock = clock; // @[:@44197.4]
  assign storeQ_reset = reset; // @[:@44198.4]
  assign storeQ_io_bbStart = GA_io_bbStart; // @[LSQAXI.scala 210:21:@44543.4]
  assign storeQ_io_bbStoreOffsets_0 = GA_io_bbStoreOffsets_0; // @[LSQAXI.scala 211:28:@44544.4]
  assign storeQ_io_bbStoreOffsets_1 = GA_io_bbStoreOffsets_1; // @[LSQAXI.scala 211:28:@44545.4]
  assign storeQ_io_bbStoreOffsets_2 = GA_io_bbStoreOffsets_2; // @[LSQAXI.scala 211:28:@44546.4]
  assign storeQ_io_bbStoreOffsets_3 = GA_io_bbStoreOffsets_3; // @[LSQAXI.scala 211:28:@44547.4]
  assign storeQ_io_bbStoreOffsets_4 = GA_io_bbStoreOffsets_4; // @[LSQAXI.scala 211:28:@44548.4]
  assign storeQ_io_bbStoreOffsets_5 = GA_io_bbStoreOffsets_5; // @[LSQAXI.scala 211:28:@44549.4]
  assign storeQ_io_bbStoreOffsets_6 = GA_io_bbStoreOffsets_6; // @[LSQAXI.scala 211:28:@44550.4]
  assign storeQ_io_bbStoreOffsets_7 = GA_io_bbStoreOffsets_7; // @[LSQAXI.scala 211:28:@44551.4]
  assign storeQ_io_bbStoreOffsets_8 = GA_io_bbStoreOffsets_8; // @[LSQAXI.scala 211:28:@44552.4]
  assign storeQ_io_bbStoreOffsets_9 = GA_io_bbStoreOffsets_9; // @[LSQAXI.scala 211:28:@44553.4]
  assign storeQ_io_bbStoreOffsets_10 = GA_io_bbStoreOffsets_10; // @[LSQAXI.scala 211:28:@44554.4]
  assign storeQ_io_bbStoreOffsets_11 = GA_io_bbStoreOffsets_11; // @[LSQAXI.scala 211:28:@44555.4]
  assign storeQ_io_bbStoreOffsets_12 = GA_io_bbStoreOffsets_12; // @[LSQAXI.scala 211:28:@44556.4]
  assign storeQ_io_bbStoreOffsets_13 = GA_io_bbStoreOffsets_13; // @[LSQAXI.scala 211:28:@44557.4]
  assign storeQ_io_bbStoreOffsets_14 = GA_io_bbStoreOffsets_14; // @[LSQAXI.scala 211:28:@44558.4]
  assign storeQ_io_bbStoreOffsets_15 = GA_io_bbStoreOffsets_15; // @[LSQAXI.scala 211:28:@44559.4]
  assign storeQ_io_bbNumStores = GA_io_bbNumStores; // @[LSQAXI.scala 213:25:@44576.4]
  assign storeQ_io_loadTail = loadTail[3:0]; // @[LSQAXI.scala 204:22:@44492.4]
  assign storeQ_io_loadHead = loadHead[3:0]; // @[LSQAXI.scala 205:22:@44493.4]
  assign storeQ_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQAXI.scala 206:23:@44494.4]
  assign storeQ_io_loadAddressDone_0 = loadQ_io_loadAddrDone_0; // @[LSQAXI.scala 207:29:@44495.4]
  assign storeQ_io_loadAddressDone_1 = loadQ_io_loadAddrDone_1; // @[LSQAXI.scala 207:29:@44496.4]
  assign storeQ_io_loadAddressDone_2 = loadQ_io_loadAddrDone_2; // @[LSQAXI.scala 207:29:@44497.4]
  assign storeQ_io_loadAddressDone_3 = loadQ_io_loadAddrDone_3; // @[LSQAXI.scala 207:29:@44498.4]
  assign storeQ_io_loadAddressDone_4 = loadQ_io_loadAddrDone_4; // @[LSQAXI.scala 207:29:@44499.4]
  assign storeQ_io_loadAddressDone_5 = loadQ_io_loadAddrDone_5; // @[LSQAXI.scala 207:29:@44500.4]
  assign storeQ_io_loadAddressDone_6 = loadQ_io_loadAddrDone_6; // @[LSQAXI.scala 207:29:@44501.4]
  assign storeQ_io_loadAddressDone_7 = loadQ_io_loadAddrDone_7; // @[LSQAXI.scala 207:29:@44502.4]
  assign storeQ_io_loadAddressDone_8 = loadQ_io_loadAddrDone_8; // @[LSQAXI.scala 207:29:@44503.4]
  assign storeQ_io_loadAddressDone_9 = loadQ_io_loadAddrDone_9; // @[LSQAXI.scala 207:29:@44504.4]
  assign storeQ_io_loadAddressDone_10 = loadQ_io_loadAddrDone_10; // @[LSQAXI.scala 207:29:@44505.4]
  assign storeQ_io_loadAddressDone_11 = loadQ_io_loadAddrDone_11; // @[LSQAXI.scala 207:29:@44506.4]
  assign storeQ_io_loadAddressDone_12 = loadQ_io_loadAddrDone_12; // @[LSQAXI.scala 207:29:@44507.4]
  assign storeQ_io_loadAddressDone_13 = loadQ_io_loadAddrDone_13; // @[LSQAXI.scala 207:29:@44508.4]
  assign storeQ_io_loadAddressDone_14 = loadQ_io_loadAddrDone_14; // @[LSQAXI.scala 207:29:@44509.4]
  assign storeQ_io_loadAddressDone_15 = loadQ_io_loadAddrDone_15; // @[LSQAXI.scala 207:29:@44510.4]
  assign storeQ_io_loadDataDone_0 = loadQ_io_loadDataDone_0; // @[LSQAXI.scala 208:26:@44511.4]
  assign storeQ_io_loadDataDone_1 = loadQ_io_loadDataDone_1; // @[LSQAXI.scala 208:26:@44512.4]
  assign storeQ_io_loadDataDone_2 = loadQ_io_loadDataDone_2; // @[LSQAXI.scala 208:26:@44513.4]
  assign storeQ_io_loadDataDone_3 = loadQ_io_loadDataDone_3; // @[LSQAXI.scala 208:26:@44514.4]
  assign storeQ_io_loadDataDone_4 = loadQ_io_loadDataDone_4; // @[LSQAXI.scala 208:26:@44515.4]
  assign storeQ_io_loadDataDone_5 = loadQ_io_loadDataDone_5; // @[LSQAXI.scala 208:26:@44516.4]
  assign storeQ_io_loadDataDone_6 = loadQ_io_loadDataDone_6; // @[LSQAXI.scala 208:26:@44517.4]
  assign storeQ_io_loadDataDone_7 = loadQ_io_loadDataDone_7; // @[LSQAXI.scala 208:26:@44518.4]
  assign storeQ_io_loadDataDone_8 = loadQ_io_loadDataDone_8; // @[LSQAXI.scala 208:26:@44519.4]
  assign storeQ_io_loadDataDone_9 = loadQ_io_loadDataDone_9; // @[LSQAXI.scala 208:26:@44520.4]
  assign storeQ_io_loadDataDone_10 = loadQ_io_loadDataDone_10; // @[LSQAXI.scala 208:26:@44521.4]
  assign storeQ_io_loadDataDone_11 = loadQ_io_loadDataDone_11; // @[LSQAXI.scala 208:26:@44522.4]
  assign storeQ_io_loadDataDone_12 = loadQ_io_loadDataDone_12; // @[LSQAXI.scala 208:26:@44523.4]
  assign storeQ_io_loadDataDone_13 = loadQ_io_loadDataDone_13; // @[LSQAXI.scala 208:26:@44524.4]
  assign storeQ_io_loadDataDone_14 = loadQ_io_loadDataDone_14; // @[LSQAXI.scala 208:26:@44525.4]
  assign storeQ_io_loadDataDone_15 = loadQ_io_loadDataDone_15; // @[LSQAXI.scala 208:26:@44526.4]
  assign storeQ_io_loadAddressQueue_0 = loadQ_io_loadAddrQueue_0; // @[LSQAXI.scala 209:30:@44527.4]
  assign storeQ_io_loadAddressQueue_1 = loadQ_io_loadAddrQueue_1; // @[LSQAXI.scala 209:30:@44528.4]
  assign storeQ_io_loadAddressQueue_2 = loadQ_io_loadAddrQueue_2; // @[LSQAXI.scala 209:30:@44529.4]
  assign storeQ_io_loadAddressQueue_3 = loadQ_io_loadAddrQueue_3; // @[LSQAXI.scala 209:30:@44530.4]
  assign storeQ_io_loadAddressQueue_4 = loadQ_io_loadAddrQueue_4; // @[LSQAXI.scala 209:30:@44531.4]
  assign storeQ_io_loadAddressQueue_5 = loadQ_io_loadAddrQueue_5; // @[LSQAXI.scala 209:30:@44532.4]
  assign storeQ_io_loadAddressQueue_6 = loadQ_io_loadAddrQueue_6; // @[LSQAXI.scala 209:30:@44533.4]
  assign storeQ_io_loadAddressQueue_7 = loadQ_io_loadAddrQueue_7; // @[LSQAXI.scala 209:30:@44534.4]
  assign storeQ_io_loadAddressQueue_8 = loadQ_io_loadAddrQueue_8; // @[LSQAXI.scala 209:30:@44535.4]
  assign storeQ_io_loadAddressQueue_9 = loadQ_io_loadAddrQueue_9; // @[LSQAXI.scala 209:30:@44536.4]
  assign storeQ_io_loadAddressQueue_10 = loadQ_io_loadAddrQueue_10; // @[LSQAXI.scala 209:30:@44537.4]
  assign storeQ_io_loadAddressQueue_11 = loadQ_io_loadAddrQueue_11; // @[LSQAXI.scala 209:30:@44538.4]
  assign storeQ_io_loadAddressQueue_12 = loadQ_io_loadAddrQueue_12; // @[LSQAXI.scala 209:30:@44539.4]
  assign storeQ_io_loadAddressQueue_13 = loadQ_io_loadAddrQueue_13; // @[LSQAXI.scala 209:30:@44540.4]
  assign storeQ_io_loadAddressQueue_14 = loadQ_io_loadAddrQueue_14; // @[LSQAXI.scala 209:30:@44541.4]
  assign storeQ_io_loadAddressQueue_15 = loadQ_io_loadAddrQueue_15; // @[LSQAXI.scala 209:30:@44542.4]
  assign storeQ_io_storeDataEnable_0 = STORE_DATA_PORT_LSQ_a_io_storeDataEnable; // @[LSQAXI.scala 221:29:@44644.4]
  assign storeQ_io_dataFromStorePorts_0 = STORE_DATA_PORT_LSQ_a_io_dataToStoreQueue; // @[LSQAXI.scala 222:32:@44645.4]
  assign storeQ_io_storeAddrEnable_0 = STORE_ADDR_PORT_LSQ_a_io_storeDataEnable; // @[LSQAXI.scala 223:29:@44646.4]
  assign storeQ_io_addressFromStorePorts_0 = sAddressPorts_0_addrToStoreQueue[30:0]; // @[LSQAXI.scala 224:35:@44647.4]
  assign storeQ_io_storeQIdxOut_ready = AXIWr_io_storeQIdxInToAW_ready; // @[LSQAXI.scala 230:32:@44652.4]
  assign storeQ_io_storeQIdxIn = AXIWr_io_storeQIdxOutFromAW; // @[LSQAXI.scala 231:25:@44653.4]
  assign storeQ_io_storeQIdxInValid = AXIWr_io_storeQIdxOutFromAWValid; // @[LSQAXI.scala 232:30:@44654.4]
  assign loadQ_clock = clock; // @[:@44200.4]
  assign loadQ_reset = reset; // @[:@44201.4]
  assign loadQ_io_bbStart = GA_io_bbStart; // @[LSQAXI.scala 178:20:@44395.4]
  assign loadQ_io_bbLoadOffsets_0 = GA_io_bbLoadOffsets_0; // @[LSQAXI.scala 179:26:@44396.4]
  assign loadQ_io_bbLoadOffsets_1 = GA_io_bbLoadOffsets_1; // @[LSQAXI.scala 179:26:@44397.4]
  assign loadQ_io_bbLoadOffsets_2 = GA_io_bbLoadOffsets_2; // @[LSQAXI.scala 179:26:@44398.4]
  assign loadQ_io_bbLoadOffsets_3 = GA_io_bbLoadOffsets_3; // @[LSQAXI.scala 179:26:@44399.4]
  assign loadQ_io_bbLoadOffsets_4 = GA_io_bbLoadOffsets_4; // @[LSQAXI.scala 179:26:@44400.4]
  assign loadQ_io_bbLoadOffsets_5 = GA_io_bbLoadOffsets_5; // @[LSQAXI.scala 179:26:@44401.4]
  assign loadQ_io_bbLoadOffsets_6 = GA_io_bbLoadOffsets_6; // @[LSQAXI.scala 179:26:@44402.4]
  assign loadQ_io_bbLoadOffsets_7 = GA_io_bbLoadOffsets_7; // @[LSQAXI.scala 179:26:@44403.4]
  assign loadQ_io_bbLoadOffsets_8 = GA_io_bbLoadOffsets_8; // @[LSQAXI.scala 179:26:@44404.4]
  assign loadQ_io_bbLoadOffsets_9 = GA_io_bbLoadOffsets_9; // @[LSQAXI.scala 179:26:@44405.4]
  assign loadQ_io_bbLoadOffsets_10 = GA_io_bbLoadOffsets_10; // @[LSQAXI.scala 179:26:@44406.4]
  assign loadQ_io_bbLoadOffsets_11 = GA_io_bbLoadOffsets_11; // @[LSQAXI.scala 179:26:@44407.4]
  assign loadQ_io_bbLoadOffsets_12 = GA_io_bbLoadOffsets_12; // @[LSQAXI.scala 179:26:@44408.4]
  assign loadQ_io_bbLoadOffsets_13 = GA_io_bbLoadOffsets_13; // @[LSQAXI.scala 179:26:@44409.4]
  assign loadQ_io_bbLoadOffsets_14 = GA_io_bbLoadOffsets_14; // @[LSQAXI.scala 179:26:@44410.4]
  assign loadQ_io_bbLoadOffsets_15 = GA_io_bbLoadOffsets_15; // @[LSQAXI.scala 179:26:@44411.4]
  assign loadQ_io_bbNumLoads = GA_io_bbNumLoads; // @[LSQAXI.scala 181:23:@44428.4]
  assign loadQ_io_storeTail = storeTail[3:0]; // @[LSQAXI.scala 171:22:@44328.4]
  assign loadQ_io_storeHead = storeHead[3:0]; // @[LSQAXI.scala 172:22:@44329.4]
  assign loadQ_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQAXI.scala 173:23:@44330.4]
  assign loadQ_io_storeAddrDone_0 = storeQ_io_storeAddrDone_0; // @[LSQAXI.scala 174:26:@44331.4]
  assign loadQ_io_storeAddrDone_1 = storeQ_io_storeAddrDone_1; // @[LSQAXI.scala 174:26:@44332.4]
  assign loadQ_io_storeAddrDone_2 = storeQ_io_storeAddrDone_2; // @[LSQAXI.scala 174:26:@44333.4]
  assign loadQ_io_storeAddrDone_3 = storeQ_io_storeAddrDone_3; // @[LSQAXI.scala 174:26:@44334.4]
  assign loadQ_io_storeAddrDone_4 = storeQ_io_storeAddrDone_4; // @[LSQAXI.scala 174:26:@44335.4]
  assign loadQ_io_storeAddrDone_5 = storeQ_io_storeAddrDone_5; // @[LSQAXI.scala 174:26:@44336.4]
  assign loadQ_io_storeAddrDone_6 = storeQ_io_storeAddrDone_6; // @[LSQAXI.scala 174:26:@44337.4]
  assign loadQ_io_storeAddrDone_7 = storeQ_io_storeAddrDone_7; // @[LSQAXI.scala 174:26:@44338.4]
  assign loadQ_io_storeAddrDone_8 = storeQ_io_storeAddrDone_8; // @[LSQAXI.scala 174:26:@44339.4]
  assign loadQ_io_storeAddrDone_9 = storeQ_io_storeAddrDone_9; // @[LSQAXI.scala 174:26:@44340.4]
  assign loadQ_io_storeAddrDone_10 = storeQ_io_storeAddrDone_10; // @[LSQAXI.scala 174:26:@44341.4]
  assign loadQ_io_storeAddrDone_11 = storeQ_io_storeAddrDone_11; // @[LSQAXI.scala 174:26:@44342.4]
  assign loadQ_io_storeAddrDone_12 = storeQ_io_storeAddrDone_12; // @[LSQAXI.scala 174:26:@44343.4]
  assign loadQ_io_storeAddrDone_13 = storeQ_io_storeAddrDone_13; // @[LSQAXI.scala 174:26:@44344.4]
  assign loadQ_io_storeAddrDone_14 = storeQ_io_storeAddrDone_14; // @[LSQAXI.scala 174:26:@44345.4]
  assign loadQ_io_storeAddrDone_15 = storeQ_io_storeAddrDone_15; // @[LSQAXI.scala 174:26:@44346.4]
  assign loadQ_io_storeDataDone_0 = storeQ_io_storeDataDone_0; // @[LSQAXI.scala 175:26:@44347.4]
  assign loadQ_io_storeDataDone_1 = storeQ_io_storeDataDone_1; // @[LSQAXI.scala 175:26:@44348.4]
  assign loadQ_io_storeDataDone_2 = storeQ_io_storeDataDone_2; // @[LSQAXI.scala 175:26:@44349.4]
  assign loadQ_io_storeDataDone_3 = storeQ_io_storeDataDone_3; // @[LSQAXI.scala 175:26:@44350.4]
  assign loadQ_io_storeDataDone_4 = storeQ_io_storeDataDone_4; // @[LSQAXI.scala 175:26:@44351.4]
  assign loadQ_io_storeDataDone_5 = storeQ_io_storeDataDone_5; // @[LSQAXI.scala 175:26:@44352.4]
  assign loadQ_io_storeDataDone_6 = storeQ_io_storeDataDone_6; // @[LSQAXI.scala 175:26:@44353.4]
  assign loadQ_io_storeDataDone_7 = storeQ_io_storeDataDone_7; // @[LSQAXI.scala 175:26:@44354.4]
  assign loadQ_io_storeDataDone_8 = storeQ_io_storeDataDone_8; // @[LSQAXI.scala 175:26:@44355.4]
  assign loadQ_io_storeDataDone_9 = storeQ_io_storeDataDone_9; // @[LSQAXI.scala 175:26:@44356.4]
  assign loadQ_io_storeDataDone_10 = storeQ_io_storeDataDone_10; // @[LSQAXI.scala 175:26:@44357.4]
  assign loadQ_io_storeDataDone_11 = storeQ_io_storeDataDone_11; // @[LSQAXI.scala 175:26:@44358.4]
  assign loadQ_io_storeDataDone_12 = storeQ_io_storeDataDone_12; // @[LSQAXI.scala 175:26:@44359.4]
  assign loadQ_io_storeDataDone_13 = storeQ_io_storeDataDone_13; // @[LSQAXI.scala 175:26:@44360.4]
  assign loadQ_io_storeDataDone_14 = storeQ_io_storeDataDone_14; // @[LSQAXI.scala 175:26:@44361.4]
  assign loadQ_io_storeDataDone_15 = storeQ_io_storeDataDone_15; // @[LSQAXI.scala 175:26:@44362.4]
  assign loadQ_io_storeAddrQueue_0 = storeQ_io_storeAddrQueue_0; // @[LSQAXI.scala 176:27:@44363.4]
  assign loadQ_io_storeAddrQueue_1 = storeQ_io_storeAddrQueue_1; // @[LSQAXI.scala 176:27:@44364.4]
  assign loadQ_io_storeAddrQueue_2 = storeQ_io_storeAddrQueue_2; // @[LSQAXI.scala 176:27:@44365.4]
  assign loadQ_io_storeAddrQueue_3 = storeQ_io_storeAddrQueue_3; // @[LSQAXI.scala 176:27:@44366.4]
  assign loadQ_io_storeAddrQueue_4 = storeQ_io_storeAddrQueue_4; // @[LSQAXI.scala 176:27:@44367.4]
  assign loadQ_io_storeAddrQueue_5 = storeQ_io_storeAddrQueue_5; // @[LSQAXI.scala 176:27:@44368.4]
  assign loadQ_io_storeAddrQueue_6 = storeQ_io_storeAddrQueue_6; // @[LSQAXI.scala 176:27:@44369.4]
  assign loadQ_io_storeAddrQueue_7 = storeQ_io_storeAddrQueue_7; // @[LSQAXI.scala 176:27:@44370.4]
  assign loadQ_io_storeAddrQueue_8 = storeQ_io_storeAddrQueue_8; // @[LSQAXI.scala 176:27:@44371.4]
  assign loadQ_io_storeAddrQueue_9 = storeQ_io_storeAddrQueue_9; // @[LSQAXI.scala 176:27:@44372.4]
  assign loadQ_io_storeAddrQueue_10 = storeQ_io_storeAddrQueue_10; // @[LSQAXI.scala 176:27:@44373.4]
  assign loadQ_io_storeAddrQueue_11 = storeQ_io_storeAddrQueue_11; // @[LSQAXI.scala 176:27:@44374.4]
  assign loadQ_io_storeAddrQueue_12 = storeQ_io_storeAddrQueue_12; // @[LSQAXI.scala 176:27:@44375.4]
  assign loadQ_io_storeAddrQueue_13 = storeQ_io_storeAddrQueue_13; // @[LSQAXI.scala 176:27:@44376.4]
  assign loadQ_io_storeAddrQueue_14 = storeQ_io_storeAddrQueue_14; // @[LSQAXI.scala 176:27:@44377.4]
  assign loadQ_io_storeAddrQueue_15 = storeQ_io_storeAddrQueue_15; // @[LSQAXI.scala 176:27:@44378.4]
  assign loadQ_io_storeDataQueue_0 = storeQ_io_storeDataQueue_0; // @[LSQAXI.scala 177:27:@44379.4]
  assign loadQ_io_storeDataQueue_1 = storeQ_io_storeDataQueue_1; // @[LSQAXI.scala 177:27:@44380.4]
  assign loadQ_io_storeDataQueue_2 = storeQ_io_storeDataQueue_2; // @[LSQAXI.scala 177:27:@44381.4]
  assign loadQ_io_storeDataQueue_3 = storeQ_io_storeDataQueue_3; // @[LSQAXI.scala 177:27:@44382.4]
  assign loadQ_io_storeDataQueue_4 = storeQ_io_storeDataQueue_4; // @[LSQAXI.scala 177:27:@44383.4]
  assign loadQ_io_storeDataQueue_5 = storeQ_io_storeDataQueue_5; // @[LSQAXI.scala 177:27:@44384.4]
  assign loadQ_io_storeDataQueue_6 = storeQ_io_storeDataQueue_6; // @[LSQAXI.scala 177:27:@44385.4]
  assign loadQ_io_storeDataQueue_7 = storeQ_io_storeDataQueue_7; // @[LSQAXI.scala 177:27:@44386.4]
  assign loadQ_io_storeDataQueue_8 = storeQ_io_storeDataQueue_8; // @[LSQAXI.scala 177:27:@44387.4]
  assign loadQ_io_storeDataQueue_9 = storeQ_io_storeDataQueue_9; // @[LSQAXI.scala 177:27:@44388.4]
  assign loadQ_io_storeDataQueue_10 = storeQ_io_storeDataQueue_10; // @[LSQAXI.scala 177:27:@44389.4]
  assign loadQ_io_storeDataQueue_11 = storeQ_io_storeDataQueue_11; // @[LSQAXI.scala 177:27:@44390.4]
  assign loadQ_io_storeDataQueue_12 = storeQ_io_storeDataQueue_12; // @[LSQAXI.scala 177:27:@44391.4]
  assign loadQ_io_storeDataQueue_13 = storeQ_io_storeDataQueue_13; // @[LSQAXI.scala 177:27:@44392.4]
  assign loadQ_io_storeDataQueue_14 = storeQ_io_storeDataQueue_14; // @[LSQAXI.scala 177:27:@44393.4]
  assign loadQ_io_storeDataQueue_15 = storeQ_io_storeDataQueue_15; // @[LSQAXI.scala 177:27:@44394.4]
  assign loadQ_io_loadAddrEnable_0 = LOAD_PORT_LSQ_a_io_loadAddrEnable; // @[LSQAXI.scala 192:32:@44484.4]
  assign loadQ_io_addrFromLoadPorts_0 = LOAD_PORT_LSQ_a_io_addrToLoadQueue; // @[LSQAXI.scala 191:35:@44483.4]
  assign loadQ_io_loadPorts_0_ready = LOAD_PORT_LSQ_a_io_dataFromLoadQueue_ready; // @[LSQAXI.scala 190:27:@44482.4]
  assign loadQ_io_loadDataFromMem = AXIRd_io_loadDataFromMem; // @[LSQAXI.scala 195:28:@44485.4]
  assign loadQ_io_loadQIdxForDataIn = AXIRd_io_loadQIdxForDataOut; // @[LSQAXI.scala 197:30:@44487.4]
  assign loadQ_io_loadQIdxForDataInValid = AXIRd_io_loadQIdxForDataOutValid; // @[LSQAXI.scala 198:35:@44488.4]
  assign loadQ_io_loadQIdxForAddrOut_ready = AXIRd_io_loadQIdxForAddrIn_ready; // @[LSQAXI.scala 201:37:@44491.4]
  assign GA_io_loadTail = loadTail[3:0]; // @[LSQAXI.scala 155:18:@44282.4]
  assign GA_io_loadHead = loadHead[3:0]; // @[LSQAXI.scala 156:18:@44283.4]
  assign GA_io_loadEmpty = loadQ_io_loadEmpty; // @[LSQAXI.scala 157:19:@44284.4]
  assign GA_io_storeTail = storeTail[3:0]; // @[LSQAXI.scala 161:19:@44318.4]
  assign GA_io_storeHead = storeHead[3:0]; // @[LSQAXI.scala 162:19:@44319.4]
  assign GA_io_storeEmpty = storeQ_io_storeEmpty; // @[LSQAXI.scala 163:20:@44320.4]
  assign GA_io_bbStartSignals_0 = io_bbStartSignals_0; // @[LSQAXI.scala 165:24:@44322.4]
  assign GA_io_bbStartSignals_1 = io_bbStartSignals_1; // @[LSQAXI.scala 165:24:@44323.4]
  assign AXIWr_clock = clock; // @[:@44206.4]
  assign AXIWr_reset = reset; // @[:@44207.4]
  assign AXIWr_io_storeAddrToMem = storeQ_io_storeAddrToMem; // @[LSQAXI.scala 266:27:@44680.4]
  assign AXIWr_io_storeDataToMem = storeQ_io_storeDataToMem; // @[LSQAXI.scala 267:27:@44681.4]
  assign AXIWr_io_storeQIdxInToAW_valid = storeQ_io_storeQIdxOut_valid; // @[LSQAXI.scala 269:34:@44683.4]
  assign AXIWr_io_storeQIdxInToAW_bits = storeQ_io_storeQIdxOut_bits; // @[LSQAXI.scala 268:33:@44682.4]
  assign AXIWr_io_AWREADY = io_AWREADY; // @[LSQAXI.scala 286:20:@44698.4]
  assign AXIWr_io_WREADY = io_WREADY; // @[LSQAXI.scala 293:19:@44704.4]
  assign AXIWr_io_BID = io_BID; // @[LSQAXI.scala 295:16:@44705.4]
  assign AXIWr_io_BRESP = io_BRESP; // @[LSQAXI.scala 296:18:@44706.4]
  assign AXIWr_io_BVALID = io_BVALID; // @[LSQAXI.scala 297:19:@44707.4]
  assign AXIRd_clock = clock; // @[:@44209.4]
  assign AXIRd_reset = reset; // @[:@44210.4]
  assign AXIRd_io_loadAddrToMem = loadQ_io_loadAddrToMem; // @[LSQAXI.scala 236:26:@44655.4]
  assign AXIRd_io_loadQIdxForAddrIn_valid = loadQ_io_loadQIdxForAddrOut_valid; // @[LSQAXI.scala 241:36:@44660.4]
  assign AXIRd_io_loadQIdxForAddrIn_bits = {{27'd0}, loadQ_io_loadQIdxForAddrOut_bits}; // @[LSQAXI.scala 240:35:@44659.4]
  assign AXIRd_io_ARREADY = io_ARREADY; // @[LSQAXI.scala 255:20:@44673.4]
  assign AXIRd_io_RID = io_RID; // @[LSQAXI.scala 258:16:@44674.4]
  assign AXIRd_io_RDATA = io_RDATA; // @[LSQAXI.scala 259:18:@44675.4]
  assign AXIRd_io_RRESP = io_RRESP; // @[LSQAXI.scala 260:18:@44676.4]
  assign AXIRd_io_RLAST = io_RLAST; // @[LSQAXI.scala 261:18:@44677.4]
  assign AXIRd_io_RVALID = io_RVALID; // @[LSQAXI.scala 262:19:@44678.4]
  assign LOAD_PORT_LSQ_a_clock = clock; // @[:@44212.4]
  assign LOAD_PORT_LSQ_a_reset = reset; // @[:@44213.4]
  assign LOAD_PORT_LSQ_a_io_addrFromPrev_valid = io_previousAndLoadPorts_0_valid; // @[LSQAXI.scala 137:23:@44225.4]
  assign LOAD_PORT_LSQ_a_io_addrFromPrev_bits = io_previousAndLoadPorts_0_bits; // @[LSQAXI.scala 137:23:@44224.4]
  assign LOAD_PORT_LSQ_a_io_portEnable = GA_io_loadPortsEnable_0; // @[LSQAXI.scala 137:23:@44223.4]
  assign LOAD_PORT_LSQ_a_io_dataToNext_ready = io_nextAndLoadPorts_0_ready; // @[LSQAXI.scala 137:23:@44222.4]
  assign LOAD_PORT_LSQ_a_io_dataFromLoadQueue_valid = loadQ_io_loadPorts_0_valid; // @[LSQAXI.scala 137:23:@44216.4]
  assign LOAD_PORT_LSQ_a_io_dataFromLoadQueue_bits = loadQ_io_loadPorts_0_bits; // @[LSQAXI.scala 137:23:@44215.4]
  assign STORE_DATA_PORT_LSQ_a_clock = clock; // @[:@44228.4]
  assign STORE_DATA_PORT_LSQ_a_reset = reset; // @[:@44229.4]
  assign STORE_DATA_PORT_LSQ_a_io_dataFromPrev_valid = io_previousAndStoreDataPorts_0_valid; // @[LSQAXI.scala 141:27:@44235.4]
  assign STORE_DATA_PORT_LSQ_a_io_dataFromPrev_bits = io_previousAndStoreDataPorts_0_bits; // @[LSQAXI.scala 141:27:@44234.4]
  assign STORE_DATA_PORT_LSQ_a_io_portEnable = GA_io_storePortsEnable_0; // @[LSQAXI.scala 141:27:@44233.4]
  assign STORE_ADDR_PORT_LSQ_a_clock = clock; // @[:@44238.4]
  assign STORE_ADDR_PORT_LSQ_a_reset = reset; // @[:@44239.4]
  assign STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_valid = io_previousAndStoreAddressPorts_0_valid; // @[LSQAXI.scala 145:30:@44245.4]
  assign STORE_ADDR_PORT_LSQ_a_io_dataFromPrev_bits = {{1'd0}, io_previousAndStoreAddressPorts_0_bits}; // @[LSQAXI.scala 145:30:@44244.4]
  assign STORE_ADDR_PORT_LSQ_a_io_portEnable = GA_io_storePortsEnable_0; // @[LSQAXI.scala 145:30:@44243.4]
endmodule
